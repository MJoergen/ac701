
`timescale 1ps / 1ps
module model_ap2_tst_pcie_2_1_rport_7x # (
    parameter        CFG_VEND_ID = 16'h10ee,
    parameter        CFG_DEV_ID = 16'h7124,
    parameter        UPSTREAM_FACING = "FALSE",    

    parameter        CFG_REV_ID =  8'h00,
    parameter        CFG_SUBSYS_VEND_ID = 16'h10ee,
    parameter        CFG_SUBSYS_ID = 16'h0007,

    parameter         EXT_PIPE_SIM = "FALSE",
    // PCIE_2_1 params
    parameter        REF_CLK_FREQ = 0,
    parameter        PCIE_EXT_CLK = "FALSE",
    parameter        PIPE_PIPELINE_STAGES = 0,

    parameter [11:0] AER_BASE_PTR = 12'h128,
    parameter        AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
    parameter        AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
    parameter [15:0] AER_CAP_ID = 16'h0001,
    parameter        AER_CAP_MULTIHEADER = "FALSE",
    parameter [11:0] AER_CAP_NEXTPTR = 12'h160,
    parameter        AER_CAP_ON = "FALSE",
    parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000,
    parameter        AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE",
    parameter [3:0]  AER_CAP_VERSION = 4'h1,
    parameter        ALLOW_X8_GEN2 = "FALSE",

    parameter [31:0] BAR0 = 32'hFFE00000,
    parameter [31:0] BAR1 = 32'hFFFFF800,
    parameter [31:0] BAR2 = 32'hFFFFF800,
    parameter [31:0] BAR3 = 32'h00000000,
    parameter [31:0] BAR4 = 32'h00000000,
    parameter [31:0] BAR5 = 32'h00000000,

    parameter        C_DATA_WIDTH = 64,
    parameter [7:0]  CAPABILITIES_PTR = 8'h40,
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000,
    parameter        CFG_ECRC_ERR_CPLSTAT = 0,
    parameter [23:0] CLASS_CODE = 24'h050000,
    parameter        CMD_INTX_IMPLEMENTED = "FALSE",
    parameter        CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE",
    parameter [3:0]  CPL_TIMEOUT_RANGES_SUPPORTED = 4'h2,
    parameter [6:0]  CRM_MODULE_RSTS = 7'h00,

    parameter        DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE",
    parameter        DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE",
    parameter [1:0]  DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0,
    parameter        DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE",
    parameter [1:0]  DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0,

    parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE",
    parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE",
    parameter        integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0,
    parameter        integer DEV_CAP_ENDPOINT_L1_LATENCY = 0,
    parameter        DEV_CAP_EXT_TAG_SUPPORTED = "TRUE",
    parameter        DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE",
    parameter        integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2,
    parameter        integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0,
    parameter        DEV_CAP_ROLE_BASED_ERROR = "TRUE",
    parameter        integer DEV_CAP_RSVD_14_12 = 0,
    parameter        integer DEV_CAP_RSVD_17_16 = 0,
    parameter        integer DEV_CAP_RSVD_31_29 = 0,
    parameter        DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE",
    parameter        DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE",
    parameter        DISABLE_ASPM_L1_TIMER = "FALSE",
    parameter        DISABLE_BAR_FILTERING = "FALSE",
    parameter        DISABLE_ERR_MSG = "FALSE",
    parameter        DISABLE_ID_CHECK = "FALSE",
    parameter        DISABLE_LANE_REVERSAL = "FALSE",
    parameter        DISABLE_LOCKED_FILTER = "FALSE",
    parameter        DISABLE_PPM_FILTER = "FALSE",
    parameter        DISABLE_RX_POISONED_RESP = "FALSE",
    parameter        DISABLE_RX_TC_FILTER = "FALSE",
    parameter        DISABLE_SCRAMBLING = "FALSE",
    parameter [7:0]  DNSTREAM_LINK_NUM = 8'h00,
    parameter [11:0] DSN_BASE_PTR = 12'h100,
    parameter [15:0] DSN_CAP_ID = 16'h0003,
    parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C,
    parameter        DSN_CAP_ON = "TRUE",
    parameter [3:0]  DSN_CAP_VERSION = 4'h1,
    parameter [10:0] ENABLE_MSG_ROUTE = 11'h000,
    parameter        ENABLE_RX_TD_ECRC_TRIM = "FALSE",
    parameter        ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE",
    parameter        ENTER_RVRY_EI_L0 = "TRUE",
    parameter        EXIT_LOOPBACK_ON_EI = "TRUE",
    parameter [31:0] EXPANSION_ROM = 32'hFFFFF001,
    parameter [5:0]  EXT_CFG_CAP_PTR = 6'h3F,
    parameter [9:0]  EXT_CFG_XP_CAP_PTR = 10'h3FF,
    parameter [7:0]  HEADER_TYPE = 8'h00,
    parameter [4:0]  INFER_EI = 5'h00,
    parameter [7:0]  INTERRUPT_PIN = 8'h01,
    parameter        INTERRUPT_STAT_AUTO = "TRUE",
    parameter        IS_SWITCH = "FALSE",
    parameter [9:0]  LAST_CONFIG_DWORD = 10'h3FF,
    parameter        LINK_CAP_ASPM_OPTIONALITY = "TRUE",
    parameter        integer LINK_CAP_ASPM_SUPPORT = 0,
    parameter        LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE",
    parameter        LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE",
    parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7,
    parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7,
    parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7,
    parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7,
    parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7,
    parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7,
    parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7,
    parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7,
    parameter        LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE",
    parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,
    parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,
    parameter        integer LINK_CAP_RSVD_23 = 0,
    parameter        LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE",
    parameter        EXT_PIPE_INTERFACE = "FALSE",
    parameter        integer LINK_CONTROL_RCB = 0,
    parameter        LINK_CTRL2_DEEMPHASIS = "FALSE",
    parameter        LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE",
    parameter [3:0]  LINK_CTRL2_TARGET_LINK_SPEED = 4'h2,
    parameter        LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE",
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0000,
    parameter        LL_ACK_TIMEOUT_EN = "FALSE",
    parameter        integer LL_ACK_TIMEOUT_FUNC = 0,
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000,
    parameter        LL_REPLAY_TIMEOUT_EN = "FALSE",
    parameter        integer LL_REPLAY_TIMEOUT_FUNC = 0,
    parameter [5:0]  LTSSM_MAX_LINK_WIDTH = LINK_CAP_MAX_LINK_WIDTH,
    parameter        MPS_FORCE = "FALSE",
    parameter [7:0]  MSIX_BASE_PTR = 8'h9C,
    parameter [7:0]  MSIX_CAP_ID = 8'h11,
    parameter [7:0]  MSIX_CAP_NEXTPTR = 8'h00,
    parameter        MSIX_CAP_ON = "FALSE",
    parameter        integer MSIX_CAP_PBA_BIR = 0,
    parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050,
    parameter        integer MSIX_CAP_TABLE_BIR = 0,
    parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040,
    parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000,
    parameter [7:0]  MSI_BASE_PTR = 8'h48,
    parameter        MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE",
    parameter [7:0]  MSI_CAP_ID = 8'h05,
    parameter        integer MSI_CAP_MULTIMSGCAP = 0,
    parameter        integer MSI_CAP_MULTIMSG_EXTENSION = 0,
    parameter [7:0]  MSI_CAP_NEXTPTR = 8'h60,
    parameter        MSI_CAP_ON = "FALSE",
    parameter        MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE",
    parameter        integer N_FTS_COMCLK_GEN1 = 255,
    parameter        integer N_FTS_COMCLK_GEN2 = 255,
    parameter        integer N_FTS_GEN1 = 255,
    parameter        integer N_FTS_GEN2 = 255,
    parameter [7:0]  PCIE_BASE_PTR = 8'h60,
    parameter [7:0]  PCIE_CAP_CAPABILITY_ID = 8'h10,
    parameter [3:0]  PCIE_CAP_CAPABILITY_VERSION = 4'h2,
    parameter [3:0]  PCIE_CAP_DEVICE_PORT_TYPE = 4'h0,
    parameter [7:0]  PCIE_CAP_NEXTPTR = 8'h9C,
    parameter        PCIE_CAP_ON = "TRUE",
    parameter        integer PCIE_CAP_RSVD_15_14 = 0,
    parameter        PCIE_CAP_SLOT_IMPLEMENTED = "FALSE",
    parameter        integer PCIE_REVISION = 2,
    parameter        integer PL_AUTO_CONFIG = 0,
    parameter        PL_FAST_TRAIN = "FALSE",
    parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000,
    parameter        PM_ASPML0S_TIMEOUT_EN = "FALSE",
    parameter        integer PM_ASPML0S_TIMEOUT_FUNC = 0,
    parameter        PM_ASPM_FASTEXIT = "FALSE",
    parameter [7:0]  PM_BASE_PTR = 8'h40,
    parameter        integer PM_CAP_AUXCURRENT = 0,
    parameter        PM_CAP_D1SUPPORT = "TRUE",
    parameter        PM_CAP_D2SUPPORT = "TRUE",
    parameter        PM_CAP_DSI = "FALSE",
    parameter [7:0]  PM_CAP_ID = 8'h01,
    parameter [7:0]  PM_CAP_NEXTPTR = 8'h48,
    parameter        PM_CAP_ON = "TRUE",
    parameter [4:0]  PM_CAP_PMESUPPORT = 5'h0F,
    parameter        PM_CAP_PME_CLOCK = "FALSE",
    parameter        integer PM_CAP_RSVD_04 = 0,
    parameter        integer PM_CAP_VERSION = 3,
    parameter        PM_CSR_B2B3 = "FALSE",
    parameter        PM_CSR_BPCCEN = "FALSE",
    parameter        PM_CSR_NOSOFTRST = "TRUE",
    parameter [7:0]  PM_DATA0 = 8'h01,
    parameter [7:0]  PM_DATA1 = 8'h01,
    parameter [7:0]  PM_DATA2 = 8'h01,
    parameter [7:0]  PM_DATA3 = 8'h01,
    parameter [7:0]  PM_DATA4 = 8'h01,
    parameter [7:0]  PM_DATA5 = 8'h01,
    parameter [7:0]  PM_DATA6 = 8'h01,
    parameter [7:0]  PM_DATA7 = 8'h01,
    parameter [1:0]  PM_DATA_SCALE0 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE1 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE2 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE3 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE4 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE5 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE6 = 2'h1,
    parameter [1:0]  PM_DATA_SCALE7 = 2'h1,
    parameter        PM_MF = "FALSE",
    parameter [11:0] RBAR_BASE_PTR = 12'h178,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00,
    parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00,
    parameter [15:0] RBAR_CAP_ID = 16'h0015,
    parameter [2:0]  RBAR_CAP_INDEX0 = 3'h0,
    parameter [2:0]  RBAR_CAP_INDEX1 = 3'h0,
    parameter [2:0]  RBAR_CAP_INDEX2 = 3'h0,
    parameter [2:0]  RBAR_CAP_INDEX3 = 3'h0,
    parameter [2:0]  RBAR_CAP_INDEX4 = 3'h0,
    parameter [2:0]  RBAR_CAP_INDEX5 = 3'h0,
    parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000,
    parameter        RBAR_CAP_ON = "FALSE",
    parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000,
    parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000,
    parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000,
    parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000,
    parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000,
    parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000,
    parameter [3:0]  RBAR_CAP_VERSION = 4'h1,
    parameter [2:0]  RBAR_NUM = 3'h1,
    parameter        integer RECRC_CHK = 0,
    parameter        RECRC_CHK_TRIM = "FALSE",
    parameter        REM_WIDTH = (C_DATA_WIDTH == 128) ? 2 : 1,
    parameter        ROOT_CAP_CRS_SW_VISIBILITY = "FALSE",
    parameter [1:0]  RP_AUTO_SPD = 2'h1,
    parameter [4:0]  RP_AUTO_SPD_LOOPCNT = 5'h1f,
    parameter        SELECT_DLL_IF = "FALSE",
    parameter        SIM_VERSION = "1.0",
    parameter        SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE",
    parameter        SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE",
    parameter        SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE",
    parameter        SLOT_CAP_HOTPLUG_CAPABLE = "FALSE",
    parameter        SLOT_CAP_HOTPLUG_SURPRISE = "FALSE",
    parameter        SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE",
    parameter        SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE",
    parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000,
    parameter        SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE",
    parameter        SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE",
    parameter        integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0,
    parameter [7:0]  SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00,

  parameter integer SPARE_BIT0 = 0,

    parameter        integer SPARE_BIT1 = 0,
    parameter        integer SPARE_BIT2 = 0,
    parameter        integer SPARE_BIT3 = 0,
    parameter        integer SPARE_BIT4 = 0,
    parameter        integer SPARE_BIT5 = 0,
    parameter        integer SPARE_BIT6 = 0,
    parameter        integer SPARE_BIT7 = 0,
    parameter        integer SPARE_BIT8 = 0,
    parameter [7:0]  SPARE_BYTE0 = 8'h00,
    parameter [7:0]  SPARE_BYTE1 = 8'h00,
    parameter [7:0]  SPARE_BYTE2 = 8'h00,
    parameter [7:0]  SPARE_BYTE3 = 8'h00,
    parameter [31:0] SPARE_WORD0 = 32'h00000000,
    parameter [31:0] SPARE_WORD1 = 32'h00000000,
    parameter [31:0] SPARE_WORD2 = 32'h00000000,
    parameter [31:0] SPARE_WORD3 = 32'h00000000,
    parameter        SSL_MESSAGE_AUTO = "FALSE",
    parameter        KEEP_WIDTH = C_DATA_WIDTH / 8,
    parameter        TECRC_EP_INV = "FALSE",
    parameter        TL_RBYPASS = "FALSE",
    parameter        integer TL_RX_RAM_RADDR_LATENCY = 0,
    parameter        integer TL_RX_RAM_RDATA_LATENCY = 2,
    parameter        integer TL_RX_RAM_WRITE_LATENCY = 0,
    parameter        TL_TFC_DISABLE = "FALSE",
    parameter        TL_TX_CHECKS_DISABLE = "FALSE",
    parameter        integer TL_TX_RAM_RADDR_LATENCY = 0,
    parameter        integer TL_TX_RAM_RDATA_LATENCY = 2,
    parameter        integer TL_TX_RAM_WRITE_LATENCY = 0,
    parameter        TRN_DW = "FALSE",
    parameter        TRN_NP_FC = "FALSE",
    parameter        UPCONFIG_CAPABLE = "TRUE",
    
    parameter        UR_ATOMIC = "TRUE",
    parameter        UR_CFG1 = "TRUE",
    parameter        UR_INV_REQ = "TRUE",
    parameter        UR_PRS_RESPONSE = "TRUE",
    parameter        USER_CLK2_DIV2 = "FALSE",
    parameter        integer USER_CLK_FREQ = 3,
    parameter        USE_RID_PINS = "FALSE",
    parameter        VC0_CPL_INFINITE = "TRUE",
    parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF,
    parameter        integer VC0_TOTAL_CREDITS_CD = 127,
    parameter        integer VC0_TOTAL_CREDITS_CH = 31,
    parameter        integer VC0_TOTAL_CREDITS_NPD = 24,
    parameter        integer VC0_TOTAL_CREDITS_NPH = 12,
    parameter        integer VC0_TOTAL_CREDITS_PD = 288,
    parameter        integer VC0_TOTAL_CREDITS_PH = 32,
    parameter        integer VC0_TX_LASTPACKET = 31,
    parameter [11:0] VC_BASE_PTR = 12'h10C,
    parameter [15:0] VC_CAP_ID = 16'h0002,
    parameter [11:0] VC_CAP_NEXTPTR = 12'h128,
    parameter        VC_CAP_ON = "FALSE",
    parameter        VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE",
    parameter [3:0]  VC_CAP_VERSION = 4'h1,
    parameter [11:0] VSEC_BASE_PTR = 12'h160,
    parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234,
    parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018,
    parameter [3:0]  VSEC_CAP_HDR_REVISION = 4'h1,
    parameter [15:0] VSEC_CAP_ID = 16'h000B,
    parameter        VSEC_CAP_IS_LINK_VISIBLE = "TRUE",
    parameter [11:0] VSEC_CAP_NEXTPTR = 12'h000,
    parameter        VSEC_CAP_ON = "FALSE",
    parameter [3:0]  VSEC_CAP_VERSION = 4'h1,
    parameter        PCIE_USE_MODE = "3.0",
    parameter        PCIE_GT_DEVICE = "GTX",
    parameter        PCIE_CHAN_BOND = 0,
    parameter        PCIE_PLL_SEL   = "CPLL",
    parameter        PCIE_ASYNC_EN  = "FALSE",
    parameter        PCIE_TXBUF_EN  = "FALSE"
)
(

  //----------------------------------------------------------------------------------------------------------------//
  // 1. PCI Express (pci_exp) Interface                                                                             //
  //----------------------------------------------------------------------------------------------------------------//

  // Tx
  output [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pci_exp_txn,
  output [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pci_exp_txp,

  // Rx
  input  [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pci_exp_rxn,
  input  [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pci_exp_rxp,

  //----------------------------------------------------------------------------------------------------------------//
  // 2. Clock Inputs                                                                                                //
  //----------------------------------------------------------------------------------------------------------------//
  input                                      pipe_pclk_in,
  input                                      pipe_rxusrclk_in,
  input  [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pipe_rxoutclk_in,
  input                                      pipe_dclk_in,
  input                                      pipe_userclk1_in,
  input                                      pipe_userclk2_in,
  input                                      pipe_oobclk_in,
  input                                      pipe_mmcm_lock_in,

  output                                     pipe_txoutclk_out,
  output [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pipe_rxoutclk_out,
  output [(LINK_CAP_MAX_LINK_WIDTH - 1) : 0] pipe_pclk_sel_out,
  output                                     pipe_gen3_out,

  //----------------------------------------------------------------------------------------------------------------//
  // 3. AXI-S Interface                                                                                             //
  //----------------------------------------------------------------------------------------------------------------//

  // Common
  output                                     user_clk_out,
  output reg                                 user_reset_out,
  output reg                                 user_lnk_up,

  // AXI TX
  //-----------
  output  [5:0]                              tx_buf_av,
  output                                     tx_err_drop,
  output                                     tx_cfg_req,
  input  [C_DATA_WIDTH-1:0]                  s_axis_tx_tdata,
  input                                      s_axis_tx_tvalid,
  output                                     s_axis_tx_tready,
  input    [KEEP_WIDTH-1:0]                  s_axis_tx_tkeep,
  input                                      s_axis_tx_tlast,
  input               [3:0]                  s_axis_tx_tuser,
  input                                      tx_cfg_gnt,

  // AXI RX
  //-----------
  output [C_DATA_WIDTH-1:0]                  m_axis_rx_tdata,
  output                                     m_axis_rx_tvalid,
  input                                      m_axis_rx_tready,
  output   [KEEP_WIDTH-1:0]                  m_axis_rx_tkeep,
  output                                     m_axis_rx_tlast,
  output             [21:0]                  m_axis_rx_tuser,
  input                                      rx_np_ok,
  input                                      rx_np_req,

  // Flow Control
  output  [11:0]                             fc_cpld,
  output  [7:0]                              fc_cplh,
  output  [11:0]                             fc_npd,
  output  [7:0]                              fc_nph,
  output  [11:0]                             fc_pd,
  output  [7:0]                              fc_ph,
  input   [2:0]                              fc_sel,


  //----------------------------------------------------------------------------------------------------------------//
  // 4. Configuration (CFG) Interface                                                                               //
  //----------------------------------------------------------------------------------------------------------------//

  //------------------------------------------------//
  // EP and RP                                      //
  //------------------------------------------------//
  output wire  [31:0]  cfg_mgmt_do,
  output wire          cfg_mgmt_rd_wr_done,

  output wire  [15:0]  cfg_status,
  output wire  [15:0]  cfg_command,
  output wire  [15:0]  cfg_dstatus,
  output wire  [15:0]  cfg_dcommand,
  output wire  [15:0]  cfg_lstatus,
  output wire  [15:0]  cfg_lcommand,
  output wire  [15:0]  cfg_dcommand2,
  output       [2:0]   cfg_pcie_link_state,

  output wire          cfg_pmcsr_pme_en,
  output wire  [1:0]   cfg_pmcsr_powerstate,
  output wire          cfg_pmcsr_pme_status,
  output wire          cfg_received_func_lvl_rst,

  // Management Interface
  input wire   [31:0]  cfg_mgmt_di,
  input wire   [3:0]   cfg_mgmt_byte_en,
  input wire   [9:0]   cfg_mgmt_dwaddr,
  input wire           cfg_mgmt_wr_en,
  input wire           cfg_mgmt_rd_en,
  input wire           cfg_mgmt_wr_readonly,

  // Error Reporting Interface
  input wire           cfg_err_ecrc,
  input wire           cfg_err_ur,
  input wire           cfg_err_cpl_timeout,
  input wire           cfg_err_cpl_unexpect,
  input wire           cfg_err_cpl_abort,
  input wire           cfg_err_posted,
  input wire           cfg_err_cor,
  input wire           cfg_err_atomic_egress_blocked,
  input wire           cfg_err_internal_cor,
  input wire           cfg_err_malformed,
  input wire           cfg_err_mc_blocked,
  input wire           cfg_err_poisoned,
  input wire           cfg_err_norecovery,
  input wire  [47:0]   cfg_err_tlp_cpl_header,
  output wire          cfg_err_cpl_rdy,
  input wire           cfg_err_locked,
  input wire           cfg_err_acs,
  input wire           cfg_err_internal_uncor,

  input wire           cfg_trn_pending,
  input wire           cfg_pm_halt_aspm_l0s,
  input wire           cfg_pm_halt_aspm_l1,
  input wire           cfg_pm_force_state_en,
  input wire   [1:0]   cfg_pm_force_state,

  input wire  [63:0]   cfg_dsn,
  output               cfg_msg_received,
  output      [15:0]   cfg_msg_data,

  //------------------------------------------------//
  // EP Only                                        //
  //------------------------------------------------//

  // Interrupt Interface Signals
  input wire           cfg_interrupt,
  output wire          cfg_interrupt_rdy,
  input wire           cfg_interrupt_assert,
  input wire   [7:0]   cfg_interrupt_di,
  output wire  [7:0]   cfg_interrupt_do,
  output wire  [2:0]   cfg_interrupt_mmenable,
  output wire          cfg_interrupt_msienable,
  output wire          cfg_interrupt_msixenable,
  output wire          cfg_interrupt_msixfm,
  input wire           cfg_interrupt_stat,
  input wire   [4:0]   cfg_pciecap_interrupt_msgnum,


  output               cfg_to_turnoff,
  input wire           cfg_turnoff_ok,
  output wire  [7:0]   cfg_bus_number,
  output wire  [4:0]   cfg_device_number,
  output wire  [2:0]   cfg_function_number,
  input wire           cfg_pm_wake,

  output wire          cfg_msg_received_pm_as_nak,
  output wire          cfg_msg_received_setslotpowerlimit,

  //------------------------------------------------//
  // RP Only                                        //
  //------------------------------------------------//
  input wire           cfg_pm_send_pme_to,
  input  wire  [7:0]   cfg_ds_bus_number,
  input  wire  [4:0]   cfg_ds_device_number,
  input  wire  [2:0]   cfg_ds_function_number,

  input wire           cfg_mgmt_wr_rw1c_as_rw,

  output wire          cfg_bridge_serr_en,
  output wire          cfg_slot_control_electromech_il_ctl_pulse,
  output wire          cfg_root_control_syserr_corr_err_en,
  output wire          cfg_root_control_syserr_non_fatal_err_en,
  output wire          cfg_root_control_syserr_fatal_err_en,
  output wire          cfg_root_control_pme_int_en,
  output wire          cfg_aer_rooterr_corr_err_reporting_en,
  output wire          cfg_aer_rooterr_non_fatal_err_reporting_en,
  output wire          cfg_aer_rooterr_fatal_err_reporting_en,
  output wire          cfg_aer_rooterr_corr_err_received,
  output wire          cfg_aer_rooterr_non_fatal_err_received,
  output wire          cfg_aer_rooterr_fatal_err_received,

  output wire          cfg_msg_received_err_cor,
  output wire          cfg_msg_received_err_non_fatal,
  output wire          cfg_msg_received_err_fatal,
  output wire          cfg_msg_received_pm_pme,
  output wire          cfg_msg_received_pme_to_ack,
  output wire          cfg_msg_received_assert_int_a,
  output wire          cfg_msg_received_assert_int_b,
  output wire          cfg_msg_received_assert_int_c,
  output wire          cfg_msg_received_assert_int_d,
  output wire          cfg_msg_received_deassert_int_a,
  output wire          cfg_msg_received_deassert_int_b,
  output wire          cfg_msg_received_deassert_int_c,
  output wire          cfg_msg_received_deassert_int_d,
  //----------------------------------------------------------------------------------------------------------------//
  // 5. Physical Layer Control and Status (PL) Interface                                                            //
  //----------------------------------------------------------------------------------------------------------------//

  //------------------------------------------------//
  // EP and RP                                      //
  //------------------------------------------------//
  input wire   [1:0]   pl_directed_link_change,
  input wire   [1:0]   pl_directed_link_width,
  input wire           pl_directed_link_speed,
  input wire           pl_directed_link_auton,
  input wire           pl_upstream_prefer_deemph,



  output wire          pl_sel_lnk_rate,
  output wire  [1:0]   pl_sel_lnk_width,
  output wire  [5:0]   pl_ltssm_state,
  output wire  [1:0]   pl_lane_reversal_mode,

  output wire          pl_phy_lnk_up,
  output wire  [2:0]   pl_tx_pm_state,
  output wire  [1:0]   pl_rx_pm_state,

  output wire          pl_link_upcfg_cap,
  output wire          pl_link_gen2_cap,
  output wire          pl_link_partner_gen2_supported,
  output wire  [2:0]   pl_initial_link_width,

  output wire          pl_directed_change_done,

  //------------------------------------------------//
  // EP Only                                        //
  //------------------------------------------------//
  output wire          pl_received_hot_rst,

  //------------------------------------------------//
  // RP Only                                        //
  //------------------------------------------------//
  input wire           pl_transmit_hot_rst,
  input wire           pl_downstream_deemph_source,

  //----------------------------------------------------------------------------------------------------------------//
  // 6. AER interface                                                                                               //
  //----------------------------------------------------------------------------------------------------------------//

  input wire [127:0]   cfg_err_aer_headerlog,
  input wire   [4:0]   cfg_aer_interrupt_msgnum,
  output wire          cfg_err_aer_headerlog_set,
  output wire          cfg_aer_ecrc_check_en,
  output wire          cfg_aer_ecrc_gen_en,

  //----------------------------------------------------------------------------------------------------------------//
  // 7. VC interface                                                                                                //
  //----------------------------------------------------------------------------------------------------------------//

  output wire [6:0]    cfg_vc_tcvc_map,

  //----------------------------------------------------------------------------------------------------------------//
  // PIPE PORTS to TOP Level For PIPE SIMULATION with 3rd Party IP/BFM/Xilinx BFM
  //----------------------------------------------------------------------------------------------------------------//
  input wire   [11:0]  common_commands_in,
  input wire   [24:0]  pipe_rx_0_sigs,
  input wire   [24:0]  pipe_rx_1_sigs,
  input wire   [24:0]  pipe_rx_2_sigs,
  input wire   [24:0]  pipe_rx_3_sigs,
  input wire   [24:0]  pipe_rx_4_sigs,
  input wire   [24:0]  pipe_rx_5_sigs,
  input wire   [24:0]  pipe_rx_6_sigs,
  input wire   [24:0]  pipe_rx_7_sigs,

  output wire  [11:0]  common_commands_out,
  output wire  [24:0]  pipe_tx_0_sigs,
  output wire  [24:0]  pipe_tx_1_sigs,
  output wire  [24:0]  pipe_tx_2_sigs,
  output wire  [24:0]  pipe_tx_3_sigs,
  output wire  [24:0]  pipe_tx_4_sigs,
  output wire  [24:0]  pipe_tx_5_sigs,
  output wire  [24:0]  pipe_tx_6_sigs,
  output wire  [24:0]  pipe_tx_7_sigs,
  //----------------------------------------------------------------------------------------------------------------//
  // 8. System(SYS) Interface                                                                                       //
  //----------------------------------------------------------------------------------------------------------------//

  input wire           pipe_mmcm_rst_n,        // Async      | Async
  input wire           sys_clk,
  input wire           sys_rst_n
);

  wire                 user_clk;
  wire                 user_clk2;
  wire                 pipe_clk;

  wire [15:0]          cfg_vend_id        = CFG_VEND_ID;
  wire [15:0]          cfg_dev_id         = CFG_DEV_ID;
  wire [7:0]           cfg_rev_id         = CFG_REV_ID;
  wire [15:0]          cfg_subsys_vend_id = CFG_SUBSYS_VEND_ID;
  wire [15:0]          cfg_subsys_id      = CFG_SUBSYS_ID;

  // PIPE Interface Wires
  wire                 phy_rdy_n;
  wire                 pipe_rx0_polarity_gt;
  wire                 pipe_rx1_polarity_gt;
  wire                 pipe_rx2_polarity_gt;
  wire                 pipe_rx3_polarity_gt;
  wire                 pipe_rx4_polarity_gt;
  wire                 pipe_rx5_polarity_gt;
  wire                 pipe_rx6_polarity_gt;
  wire                 pipe_rx7_polarity_gt;
  wire                 pipe_tx_deemph_gt;
  wire [2:0]           pipe_tx_margin_gt;
  wire                 pipe_tx_rate_gt;
  wire                 pipe_tx_rcvr_det_gt;
  wire [1:0]           pipe_tx0_char_is_k_gt;
  wire                 pipe_tx0_compliance_gt;
  wire [15:0]          pipe_tx0_data_gt;
  wire                 pipe_tx0_elec_idle_gt;
  wire [1:0]           pipe_tx0_powerdown_gt;
  wire [1:0]           pipe_tx1_char_is_k_gt;
  wire                 pipe_tx1_compliance_gt;
  wire [15:0]          pipe_tx1_data_gt;
  wire                 pipe_tx1_elec_idle_gt;
  wire [1:0]           pipe_tx1_powerdown_gt;
  wire [1:0]           pipe_tx2_char_is_k_gt;
  wire                 pipe_tx2_compliance_gt;
  wire [15:0]          pipe_tx2_data_gt;
  wire                 pipe_tx2_elec_idle_gt;
  wire [1:0]           pipe_tx2_powerdown_gt;
  wire [1:0]           pipe_tx3_char_is_k_gt;
  wire                 pipe_tx3_compliance_gt;
  wire [15:0]          pipe_tx3_data_gt;
  wire                 pipe_tx3_elec_idle_gt;
  wire [1:0]           pipe_tx3_powerdown_gt;
  wire [1:0]           pipe_tx4_char_is_k_gt;
  wire                 pipe_tx4_compliance_gt;
  wire [15:0]          pipe_tx4_data_gt;
  wire                 pipe_tx4_elec_idle_gt;
  wire [1:0]           pipe_tx4_powerdown_gt;
  wire [1:0]           pipe_tx5_char_is_k_gt;
  wire                 pipe_tx5_compliance_gt;
  wire [15:0]          pipe_tx5_data_gt;
  wire                 pipe_tx5_elec_idle_gt;
  wire [1:0]           pipe_tx5_powerdown_gt;
  wire [1:0]           pipe_tx6_char_is_k_gt;
  wire                 pipe_tx6_compliance_gt;
  wire [15:0]          pipe_tx6_data_gt;
  wire                 pipe_tx6_elec_idle_gt;
  wire [1:0]           pipe_tx6_powerdown_gt;
  wire [1:0]           pipe_tx7_char_is_k_gt;
  wire                 pipe_tx7_compliance_gt;
  wire [15:0]          pipe_tx7_data_gt;
  wire                 pipe_tx7_elec_idle_gt;
  wire [1:0]           pipe_tx7_powerdown_gt;

  wire                 pipe_rx0_chanisaligned_gt;
  wire  [1:0]          pipe_rx0_char_is_k_gt;
  wire  [15:0]         pipe_rx0_data_gt;
  wire                 pipe_rx0_elec_idle_gt;
  wire                 pipe_rx0_phy_status_gt;
  wire  [2:0]          pipe_rx0_status_gt;
  wire                 pipe_rx0_valid_gt;
  wire                 pipe_rx1_chanisaligned_gt;
  wire  [1:0]          pipe_rx1_char_is_k_gt;
  wire  [15:0]         pipe_rx1_data_gt;
  wire                 pipe_rx1_elec_idle_gt;
  wire                 pipe_rx1_phy_status_gt;
  wire  [2:0]          pipe_rx1_status_gt;
  wire                 pipe_rx1_valid_gt;
  wire                 pipe_rx2_chanisaligned_gt;
  wire  [1:0]          pipe_rx2_char_is_k_gt;
  wire  [15:0]         pipe_rx2_data_gt;
  wire                 pipe_rx2_elec_idle_gt;
  wire                 pipe_rx2_phy_status_gt;
  wire  [2:0]          pipe_rx2_status_gt;
  wire                 pipe_rx2_valid_gt;
  wire                 pipe_rx3_chanisaligned_gt;
  wire  [1:0]          pipe_rx3_char_is_k_gt;
  wire  [15:0]         pipe_rx3_data_gt;
  wire                 pipe_rx3_elec_idle_gt;
  wire                 pipe_rx3_phy_status_gt;
  wire  [2:0]          pipe_rx3_status_gt;
  wire                 pipe_rx3_valid_gt;
  wire                 pipe_rx4_chanisaligned_gt;
  wire  [1:0]          pipe_rx4_char_is_k_gt;
  wire  [15:0]         pipe_rx4_data_gt;
  wire                 pipe_rx4_elec_idle_gt;
  wire                 pipe_rx4_phy_status_gt;
  wire  [2:0]          pipe_rx4_status_gt;
  wire                 pipe_rx4_valid_gt;
  wire                 pipe_rx5_chanisaligned_gt;
  wire  [1:0]          pipe_rx5_char_is_k_gt;
  wire  [15:0]         pipe_rx5_data_gt;
  wire                 pipe_rx5_elec_idle_gt;
  wire                 pipe_rx5_phy_status_gt;
  wire  [2:0]          pipe_rx5_status_gt;
  wire                 pipe_rx5_valid_gt;
  wire                 pipe_rx6_chanisaligned_gt;
  wire  [1:0]          pipe_rx6_char_is_k_gt;
  wire  [15:0]         pipe_rx6_data_gt;
  wire                 pipe_rx6_elec_idle_gt;
  wire                 pipe_rx6_phy_status_gt;
  wire  [2:0]          pipe_rx6_status_gt;
  wire                 pipe_rx6_valid_gt;
  wire                 pipe_rx7_chanisaligned_gt;
  wire  [1:0]          pipe_rx7_char_is_k_gt;
  wire  [15:0]         pipe_rx7_data_gt;
  wire                 pipe_rx7_elec_idle_gt;
  wire                 pipe_rx7_phy_status_gt;
  wire  [2:0]          pipe_rx7_status_gt;
  wire                 pipe_rx7_valid_gt;

  reg                  user_lnk_up_int;
  reg                  user_reset_int;
  reg                  bridge_reset_int;
  reg                  bridge_reset_d;
  wire                 user_rst_n;
  reg                  pl_received_hot_rst_q;
  wire                 pl_received_hot_rst_wire;
  reg                  pl_phy_lnk_up_q;
  wire                 pl_phy_lnk_up_wire;
  wire                 sys_or_hot_rst;
  wire                 trn_lnk_up;

  wire [5:0]           pl_ltssm_state_int;

  wire                 qpll_qplld;
  wire                 qpll_drp_clk;
  wire                 qpll_drp_rst_n;
  wire                 qpll_drp_ovrd; 
  wire                 qpll_drp_gen3;
  wire                 qpll_drp_start;
  wire                 pipe_rst_idle;
  wire                 pipe_qrst_idle;
  wire                 pipe_rate_idle;

  localparam        TCQ = 100;


  // Assign outputs
  assign pl_ltssm_state = pl_ltssm_state_int;
  assign pl_received_hot_rst = pl_received_hot_rst_q;
  assign pl_phy_lnk_up = pl_phy_lnk_up_q;

  // Register block outputs pl_received_hot_rst and phy_lnk_up to ease timing on block output
  assign sys_or_hot_rst = !sys_rst_n || ((UPSTREAM_FACING == "TRUE") && pl_received_hot_rst_q);
  always @(posedge user_clk_out)
  begin
    if (!sys_rst_n) begin
      pl_received_hot_rst_q <= #TCQ 1'b0;
      pl_phy_lnk_up_q       <= #TCQ 1'b0;
    end else begin
      pl_received_hot_rst_q <= #TCQ pl_received_hot_rst_wire;
      pl_phy_lnk_up_q       <= #TCQ pl_phy_lnk_up_wire;
    end
  end
  //------------------------------------------------------------------------------------------------------------------//
  // Convert incoming reset from AXI required active High                                                             //
  // to active low as that is what is required by GT and PCIe Block                                                   //
  //------------------------------------------------------------------------------------------------------------------//
  // assign sys_rst_n = ~sys_reset;

  // Generate user_lnk_up
  always @(posedge user_clk_out)
  begin
    if (!sys_rst_n) begin
      user_lnk_up <= #TCQ 1'b0;
    end else begin
      user_lnk_up <= #TCQ user_lnk_up_int;
    end
  end

  always @(posedge user_clk_out)
  begin
    if (!sys_rst_n) begin
      user_lnk_up_int <= #TCQ 1'b0;
    end else begin
      user_lnk_up_int <= #TCQ trn_lnk_up;
    end
  end

  // Generate user_reset_out                                                                                          //
  // Once user reset output of PCIE and Phy Layer is active, de-assert reset                                          //
  // Only assert reset if system reset or hot reset is seen.  Keep AXI backend/user application alive otherwise       //
  //------------------------------------------------------------------------------------------------------------------//
  always @(posedge user_clk_out or posedge sys_or_hot_rst)
  begin
    if (sys_or_hot_rst) begin
      user_reset_int <= #TCQ 1'b1;
    end else if (user_rst_n && pl_phy_lnk_up_q) begin
      user_reset_int <= #TCQ 1'b0;
    end
  end

  // Invert active low reset to active high AXI reset
  always @(posedge user_clk_out or posedge sys_or_hot_rst)
  begin
    if (sys_or_hot_rst) begin
      user_reset_out <= #TCQ 1'b1;
    end else begin
      user_reset_out <= #TCQ user_reset_int;
    end
  end

  always @(posedge user_clk_out or posedge sys_or_hot_rst)
  begin
    if (sys_or_hot_rst) begin
      bridge_reset_int <= #TCQ 1'b1;
    end else if (user_rst_n && pl_phy_lnk_up_q) begin
      bridge_reset_int <= #TCQ 1'b0;
    end
  end

  // Invert active low reset to active high AXI reset
  always @(posedge user_clk_out or posedge sys_or_hot_rst)
  begin
    if (sys_or_hot_rst) begin
      bridge_reset_d <= #TCQ 1'b1;
    end else begin
      bridge_reset_d <= #TCQ bridge_reset_int;
    end
  end

generate if (EXT_PIPE_SIM == "FALSE")
begin
  //------------------------------------------------------------------------------------------------------------------//
  // **** PCI Express Core Wrapper ****                                                                               //
  // The PCI Express Core Wrapper includes the following:                                                             //
  //   1) AXI Streaming Bridge                                                                                        //
  //   2) PCIE 2_1 Hard Block                                                                                         //
  //   3) PCIE PIPE Interface Pipeline                                                                                //
  //------------------------------------------------------------------------------------------------------------------//
model_ap2_tst_pcie_top # (
    .PIPE_PIPELINE_STAGES                     ( PIPE_PIPELINE_STAGES ),
    .AER_BASE_PTR                             ( AER_BASE_PTR ),
    .AER_CAP_ECRC_CHECK_CAPABLE               ( AER_CAP_ECRC_CHECK_CAPABLE ),
    .AER_CAP_ECRC_GEN_CAPABLE                 ( AER_CAP_ECRC_GEN_CAPABLE ),
    .AER_CAP_ID                               ( AER_CAP_ID ),
    .AER_CAP_MULTIHEADER                      ( AER_CAP_MULTIHEADER ),
    .AER_CAP_NEXTPTR                          ( AER_CAP_NEXTPTR ),
    .AER_CAP_ON                               ( AER_CAP_ON ),
    .AER_CAP_OPTIONAL_ERR_SUPPORT             ( AER_CAP_OPTIONAL_ERR_SUPPORT ),
    .AER_CAP_PERMIT_ROOTERR_UPDATE            ( AER_CAP_PERMIT_ROOTERR_UPDATE ),
    .AER_CAP_VERSION                          ( AER_CAP_VERSION ),
    .ALLOW_X8_GEN2                            ( ALLOW_X8_GEN2 ),
    .BAR0                                     ( BAR0 ),
    .BAR1                                     ( BAR1 ),
    .BAR2                                     ( BAR2 ),
    .BAR3                                     ( BAR3 ),
    .BAR4                                     ( BAR4 ),
    .BAR5                                     ( BAR5 ),
    .C_DATA_WIDTH                             ( C_DATA_WIDTH ),
    .CAPABILITIES_PTR                         ( CAPABILITIES_PTR ),
    .CARDBUS_CIS_POINTER                      ( CARDBUS_CIS_POINTER ),
    .CFG_ECRC_ERR_CPLSTAT                     ( CFG_ECRC_ERR_CPLSTAT ),
    .CLASS_CODE                               ( CLASS_CODE ),
    .CMD_INTX_IMPLEMENTED                     ( CMD_INTX_IMPLEMENTED ),
    .CPL_TIMEOUT_DISABLE_SUPPORTED            ( CPL_TIMEOUT_DISABLE_SUPPORTED ),
    .CPL_TIMEOUT_RANGES_SUPPORTED             ( CPL_TIMEOUT_RANGES_SUPPORTED ),
    .CRM_MODULE_RSTS                          ( CRM_MODULE_RSTS ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE ),
    .DEV_CAP_ENDPOINT_L0S_LATENCY             ( DEV_CAP_ENDPOINT_L0S_LATENCY ),
    .DEV_CAP_ENDPOINT_L1_LATENCY              ( DEV_CAP_ENDPOINT_L1_LATENCY ),
    .DEV_CAP_EXT_TAG_SUPPORTED                ( DEV_CAP_EXT_TAG_SUPPORTED ),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     ( DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE ),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED            ( DEV_CAP_MAX_PAYLOAD_SUPPORTED ),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        ( DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT ),
    .DEV_CAP_ROLE_BASED_ERROR                 ( DEV_CAP_ROLE_BASED_ERROR ),
    .DEV_CAP_RSVD_14_12                       ( DEV_CAP_RSVD_14_12 ),
    .DEV_CAP_RSVD_17_16                       ( DEV_CAP_RSVD_17_16 ),
    .DEV_CAP_RSVD_31_29                       ( DEV_CAP_RSVD_31_29 ),
    .DEV_CONTROL_AUX_POWER_SUPPORTED          ( DEV_CONTROL_AUX_POWER_SUPPORTED ),
    .DEV_CONTROL_EXT_TAG_DEFAULT              ( DEV_CONTROL_EXT_TAG_DEFAULT ),
    .DISABLE_ASPM_L1_TIMER                    ( DISABLE_ASPM_L1_TIMER ),
    .DISABLE_BAR_FILTERING                    ( DISABLE_BAR_FILTERING ),
    .DISABLE_ID_CHECK                         ( DISABLE_ID_CHECK ),
    .DISABLE_LANE_REVERSAL                    ( DISABLE_LANE_REVERSAL ),
    .DISABLE_RX_POISONED_RESP                 ( DISABLE_RX_POISONED_RESP ),
    .DISABLE_RX_TC_FILTER                     ( DISABLE_RX_TC_FILTER ),
    .DISABLE_SCRAMBLING                       ( DISABLE_SCRAMBLING ),
    .DNSTREAM_LINK_NUM                        ( DNSTREAM_LINK_NUM ),
    .DSN_BASE_PTR                             ( DSN_BASE_PTR ),
    .DSN_CAP_ID                               ( DSN_CAP_ID ),
    .DSN_CAP_NEXTPTR                          ( DSN_CAP_NEXTPTR ),
    .DSN_CAP_ON                               ( DSN_CAP_ON ),
    .DSN_CAP_VERSION                          ( DSN_CAP_VERSION ),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED        ( DEV_CAP2_ARI_FORWARDING_SUPPORTED ),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      ( DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED ),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED      ( DEV_CAP2_CAS128_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     ( DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED ),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    ( DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED ),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED         ( DEV_CAP2_LTR_MECHANISM_SUPPORTED ),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         ( DEV_CAP2_MAX_ENDEND_TLP_PREFIXES ),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      ( DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING ),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED         ( DEV_CAP2_TPH_COMPLETER_SUPPORTED ),
    .DISABLE_ERR_MSG                          ( DISABLE_ERR_MSG ),
    .DISABLE_LOCKED_FILTER                    ( DISABLE_LOCKED_FILTER ),
    .DISABLE_PPM_FILTER                       ( DISABLE_PPM_FILTER ),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   ( ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED ),
    .ENABLE_MSG_ROUTE                         ( ENABLE_MSG_ROUTE ),
    .ENABLE_RX_TD_ECRC_TRIM                   ( ENABLE_RX_TD_ECRC_TRIM ),
    .ENTER_RVRY_EI_L0                         ( ENTER_RVRY_EI_L0 ),
    .EXIT_LOOPBACK_ON_EI                      ( EXIT_LOOPBACK_ON_EI ),
    .EXPANSION_ROM                            ( EXPANSION_ROM ),
    .EXT_CFG_CAP_PTR                          ( EXT_CFG_CAP_PTR ),
    .EXT_CFG_XP_CAP_PTR                       ( EXT_CFG_XP_CAP_PTR ),
    .HEADER_TYPE                              ( HEADER_TYPE ),
    .INFER_EI                                 ( INFER_EI ),
    .INTERRUPT_PIN                            ( INTERRUPT_PIN ),
    .INTERRUPT_STAT_AUTO                      ( INTERRUPT_STAT_AUTO ),
    .IS_SWITCH                                ( IS_SWITCH ),
    .LAST_CONFIG_DWORD                        ( LAST_CONFIG_DWORD ),
    .LINK_CAP_ASPM_OPTIONALITY                ( LINK_CAP_ASPM_OPTIONALITY ),
    .LINK_CAP_ASPM_SUPPORT                    ( LINK_CAP_ASPM_SUPPORT ),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT          ( LINK_CAP_CLOCK_POWER_MANAGEMENT ),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   ( LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1           ( LINK_CAP_L0S_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2           ( LINK_CAP_L0S_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1            ( LINK_CAP_L1_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2            ( LINK_CAP_L1_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ( LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ),
    .LINK_CAP_MAX_LINK_SPEED                  ( LINK_CAP_MAX_LINK_SPEED ),
    .LINK_CAP_MAX_LINK_WIDTH                  ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_RSVD_23                         ( LINK_CAP_RSVD_23 ),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     ( LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE ),
    .LINK_CONTROL_RCB                         ( LINK_CONTROL_RCB ),
    .LINK_CTRL2_DEEMPHASIS                    ( LINK_CTRL2_DEEMPHASIS ),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   ( LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE ),
    .LINK_CTRL2_TARGET_LINK_SPEED             ( LINK_CTRL2_TARGET_LINK_SPEED ),
    .LINK_STATUS_SLOT_CLOCK_CONFIG            ( LINK_STATUS_SLOT_CLOCK_CONFIG ),
    .LL_ACK_TIMEOUT                           ( LL_ACK_TIMEOUT ),
    .LL_ACK_TIMEOUT_EN                        ( LL_ACK_TIMEOUT_EN ),
    .LL_ACK_TIMEOUT_FUNC                      ( LL_ACK_TIMEOUT_FUNC ),
    .LL_REPLAY_TIMEOUT                        ( LL_REPLAY_TIMEOUT ),
    .LL_REPLAY_TIMEOUT_EN                     ( LL_REPLAY_TIMEOUT_EN ),
    .LL_REPLAY_TIMEOUT_FUNC                   ( LL_REPLAY_TIMEOUT_FUNC ),
    .LTSSM_MAX_LINK_WIDTH                     ( LTSSM_MAX_LINK_WIDTH ),
    .MPS_FORCE                                ( MPS_FORCE),
    .MSI_BASE_PTR                             ( MSI_BASE_PTR ),
    .MSI_CAP_ID                               ( MSI_CAP_ID ),
    .MSI_CAP_MULTIMSGCAP                      ( MSI_CAP_MULTIMSGCAP ),
    .MSI_CAP_MULTIMSG_EXTENSION               ( MSI_CAP_MULTIMSG_EXTENSION ),
    .MSI_CAP_NEXTPTR                          ( MSI_CAP_NEXTPTR ),
    .MSI_CAP_ON                               ( MSI_CAP_ON ),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE       ( MSI_CAP_PER_VECTOR_MASKING_CAPABLE ),
    .MSI_CAP_64_BIT_ADDR_CAPABLE              ( MSI_CAP_64_BIT_ADDR_CAPABLE ),
    .MSIX_BASE_PTR                            ( MSIX_BASE_PTR ),
    .MSIX_CAP_ID                              ( MSIX_CAP_ID ),
    .MSIX_CAP_NEXTPTR                         ( MSIX_CAP_NEXTPTR ),
    .MSIX_CAP_ON                              ( MSIX_CAP_ON ),
    .MSIX_CAP_PBA_BIR                         ( MSIX_CAP_PBA_BIR ),
    .MSIX_CAP_PBA_OFFSET                      ( MSIX_CAP_PBA_OFFSET ),
    .MSIX_CAP_TABLE_BIR                       ( MSIX_CAP_TABLE_BIR ),
    .MSIX_CAP_TABLE_OFFSET                    ( MSIX_CAP_TABLE_OFFSET ),
    .MSIX_CAP_TABLE_SIZE                      ( MSIX_CAP_TABLE_SIZE ),
    .N_FTS_COMCLK_GEN1                        ( N_FTS_COMCLK_GEN1 ),
    .N_FTS_COMCLK_GEN2                        ( N_FTS_COMCLK_GEN2 ),
    .N_FTS_GEN1                               ( N_FTS_GEN1 ),
    .N_FTS_GEN2                               ( N_FTS_GEN2 ),
    .PCIE_BASE_PTR                            ( PCIE_BASE_PTR ),
    .PCIE_CAP_CAPABILITY_ID                   ( PCIE_CAP_CAPABILITY_ID ),
    .PCIE_CAP_CAPABILITY_VERSION              ( PCIE_CAP_CAPABILITY_VERSION ),
    .PCIE_CAP_DEVICE_PORT_TYPE                ( PCIE_CAP_DEVICE_PORT_TYPE ),
    .PCIE_CAP_NEXTPTR                         ( PCIE_CAP_NEXTPTR ),
    .PCIE_CAP_ON                              ( PCIE_CAP_ON ),
    .PCIE_CAP_RSVD_15_14                      ( PCIE_CAP_RSVD_15_14 ),
    .PCIE_CAP_SLOT_IMPLEMENTED                ( PCIE_CAP_SLOT_IMPLEMENTED ),
    .PCIE_REVISION                            ( PCIE_REVISION ),
    .PL_AUTO_CONFIG                           ( PL_AUTO_CONFIG ),
    .PL_FAST_TRAIN                            ( PL_FAST_TRAIN ),
    .PM_ASPML0S_TIMEOUT                       ( PM_ASPML0S_TIMEOUT ),
    .PM_ASPML0S_TIMEOUT_EN                    ( PM_ASPML0S_TIMEOUT_EN ),
    .PM_ASPML0S_TIMEOUT_FUNC                  ( PM_ASPML0S_TIMEOUT_FUNC ),
    .PM_ASPM_FASTEXIT                         ( PM_ASPM_FASTEXIT ),
    .PM_BASE_PTR                              ( PM_BASE_PTR ),
    .PM_CAP_AUXCURRENT                        ( PM_CAP_AUXCURRENT ),
    .PM_CAP_D1SUPPORT                         ( PM_CAP_D1SUPPORT ),
    .PM_CAP_D2SUPPORT                         ( PM_CAP_D2SUPPORT ),
    .PM_CAP_DSI                               ( PM_CAP_DSI ),
    .PM_CAP_ID                                ( PM_CAP_ID ),
    .PM_CAP_NEXTPTR                           ( PM_CAP_NEXTPTR ),
    .PM_CAP_ON                                ( PM_CAP_ON ),
    .PM_CAP_PME_CLOCK                         ( PM_CAP_PME_CLOCK ),
    .PM_CAP_PMESUPPORT                        ( PM_CAP_PMESUPPORT ),
    .PM_CAP_RSVD_04                           ( PM_CAP_RSVD_04 ),
    .PM_CAP_VERSION                           ( PM_CAP_VERSION ),
    .PM_CSR_B2B3                              ( PM_CSR_B2B3 ),
    .PM_CSR_BPCCEN                            ( PM_CSR_BPCCEN ),
    .PM_CSR_NOSOFTRST                         ( PM_CSR_NOSOFTRST ),
    .PM_DATA0                                 ( PM_DATA0 ),
    .PM_DATA1                                 ( PM_DATA1 ),
    .PM_DATA2                                 ( PM_DATA2 ),
    .PM_DATA3                                 ( PM_DATA3 ),
    .PM_DATA4                                 ( PM_DATA4 ),
    .PM_DATA5                                 ( PM_DATA5 ),
    .PM_DATA6                                 ( PM_DATA6 ),
    .PM_DATA7                                 ( PM_DATA7 ),
    .PM_DATA_SCALE0                           ( PM_DATA_SCALE0 ),
    .PM_DATA_SCALE1                           ( PM_DATA_SCALE1 ),
    .PM_DATA_SCALE2                           ( PM_DATA_SCALE2 ),
    .PM_DATA_SCALE3                           ( PM_DATA_SCALE3 ),
    .PM_DATA_SCALE4                           ( PM_DATA_SCALE4 ),
    .PM_DATA_SCALE5                           ( PM_DATA_SCALE5 ),
    .PM_DATA_SCALE6                           ( PM_DATA_SCALE6 ),
    .PM_DATA_SCALE7                           ( PM_DATA_SCALE7 ),
    .PM_MF                                    ( PM_MF ),
    .RBAR_BASE_PTR                            ( RBAR_BASE_PTR ),
    .RBAR_CAP_CONTROL_ENCODEDBAR0             ( RBAR_CAP_CONTROL_ENCODEDBAR0 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR1             ( RBAR_CAP_CONTROL_ENCODEDBAR1 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR2             ( RBAR_CAP_CONTROL_ENCODEDBAR2 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR3             ( RBAR_CAP_CONTROL_ENCODEDBAR3 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR4             ( RBAR_CAP_CONTROL_ENCODEDBAR4 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR5             ( RBAR_CAP_CONTROL_ENCODEDBAR5 ),
    .RBAR_CAP_ID                              ( RBAR_CAP_ID),
    .RBAR_CAP_INDEX0                          ( RBAR_CAP_INDEX0 ),
    .RBAR_CAP_INDEX1                          ( RBAR_CAP_INDEX1 ),
    .RBAR_CAP_INDEX2                          ( RBAR_CAP_INDEX2 ),
    .RBAR_CAP_INDEX3                          ( RBAR_CAP_INDEX3 ),
    .RBAR_CAP_INDEX4                          ( RBAR_CAP_INDEX4 ),
    .RBAR_CAP_INDEX5                          ( RBAR_CAP_INDEX5 ),
    .RBAR_CAP_NEXTPTR                         ( RBAR_CAP_NEXTPTR ),
    .RBAR_CAP_ON                              ( RBAR_CAP_ON ),
    .RBAR_CAP_SUP0                            ( RBAR_CAP_SUP0 ),
    .RBAR_CAP_SUP1                            ( RBAR_CAP_SUP1 ),
    .RBAR_CAP_SUP2                            ( RBAR_CAP_SUP2 ),
    .RBAR_CAP_SUP3                            ( RBAR_CAP_SUP3 ),
    .RBAR_CAP_SUP4                            ( RBAR_CAP_SUP4 ),
    .RBAR_CAP_SUP5                            ( RBAR_CAP_SUP5 ),
    .RBAR_CAP_VERSION                         ( RBAR_CAP_VERSION ),
    .RBAR_NUM                                 ( RBAR_NUM ),
    .RECRC_CHK                                ( RECRC_CHK ),
    .RECRC_CHK_TRIM                           ( RECRC_CHK_TRIM ),
    .ROOT_CAP_CRS_SW_VISIBILITY               ( ROOT_CAP_CRS_SW_VISIBILITY ),
    .RP_AUTO_SPD                              ( RP_AUTO_SPD ),
    .RP_AUTO_SPD_LOOPCNT                      ( RP_AUTO_SPD_LOOPCNT ),
    .SELECT_DLL_IF                            ( SELECT_DLL_IF ),
    .SLOT_CAP_ATT_BUTTON_PRESENT              ( SLOT_CAP_ATT_BUTTON_PRESENT ),
    .SLOT_CAP_ATT_INDICATOR_PRESENT           ( SLOT_CAP_ATT_INDICATOR_PRESENT ),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT          ( SLOT_CAP_ELEC_INTERLOCK_PRESENT ),
    .SLOT_CAP_HOTPLUG_CAPABLE                 ( SLOT_CAP_HOTPLUG_CAPABLE ),
    .SLOT_CAP_HOTPLUG_SURPRISE                ( SLOT_CAP_HOTPLUG_SURPRISE ),
    .SLOT_CAP_MRL_SENSOR_PRESENT              ( SLOT_CAP_MRL_SENSOR_PRESENT ),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        ( SLOT_CAP_NO_CMD_COMPLETED_SUPPORT ),
    .SLOT_CAP_PHYSICAL_SLOT_NUM               ( SLOT_CAP_PHYSICAL_SLOT_NUM ),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT        ( SLOT_CAP_POWER_CONTROLLER_PRESENT ),
    .SLOT_CAP_POWER_INDICATOR_PRESENT         ( SLOT_CAP_POWER_INDICATOR_PRESENT ),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE          ( SLOT_CAP_SLOT_POWER_LIMIT_SCALE ),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE          ( SLOT_CAP_SLOT_POWER_LIMIT_VALUE ),
    .SPARE_BIT0                               ( SPARE_BIT0 ),
    .SPARE_BIT1                               ( SPARE_BIT1 ),
    .SPARE_BIT2                               ( SPARE_BIT2 ),
    .SPARE_BIT3                               ( SPARE_BIT3 ),
    .SPARE_BIT4                               ( SPARE_BIT4 ),
    .SPARE_BIT5                               ( SPARE_BIT5 ),
    .SPARE_BIT6                               ( SPARE_BIT6 ),
    .SPARE_BIT7                               ( SPARE_BIT7 ),
    .SPARE_BIT8                               ( SPARE_BIT8 ),
    .SPARE_BYTE0                              ( SPARE_BYTE0 ),
    .SPARE_BYTE1                              ( SPARE_BYTE1 ),
    .SPARE_BYTE2                              ( SPARE_BYTE2 ),
    .SPARE_BYTE3                              ( SPARE_BYTE3 ),
    .SPARE_WORD0                              ( SPARE_WORD0 ),
    .SPARE_WORD1                              ( SPARE_WORD1 ),
    .SPARE_WORD2                              ( SPARE_WORD2 ),
    .SPARE_WORD3                              ( SPARE_WORD3 ),
    .SSL_MESSAGE_AUTO                         ( SSL_MESSAGE_AUTO ),
    .TECRC_EP_INV                             ( TECRC_EP_INV ),
    .TL_RBYPASS                               ( TL_RBYPASS ),
    .TL_RX_RAM_RADDR_LATENCY                  ( TL_RX_RAM_RADDR_LATENCY ),
    .TL_RX_RAM_RDATA_LATENCY                  ( TL_RX_RAM_RDATA_LATENCY ),
    .TL_RX_RAM_WRITE_LATENCY                  ( TL_RX_RAM_WRITE_LATENCY ),
    .TL_TFC_DISABLE                           ( TL_TFC_DISABLE ),
    .TL_TX_CHECKS_DISABLE                     ( TL_TX_CHECKS_DISABLE ),
    .TL_TX_RAM_RADDR_LATENCY                  ( TL_TX_RAM_RADDR_LATENCY ),
    .TL_TX_RAM_RDATA_LATENCY                  ( TL_TX_RAM_RDATA_LATENCY ),
    .TL_TX_RAM_WRITE_LATENCY                  ( TL_TX_RAM_WRITE_LATENCY ),
    .TRN_DW                                   ( TRN_DW ),
    .TRN_NP_FC                                ( TRN_NP_FC ),
    .UPCONFIG_CAPABLE                         ( UPCONFIG_CAPABLE ),
    .UPSTREAM_FACING                          ( UPSTREAM_FACING ),
    .UR_ATOMIC                                ( UR_ATOMIC ),
    .UR_CFG1                                  ( UR_CFG1 ),
    .UR_INV_REQ                               ( UR_INV_REQ ),
    .UR_PRS_RESPONSE                          ( UR_PRS_RESPONSE ),
    .USER_CLK2_DIV2                           ( USER_CLK2_DIV2 ),
    .USER_CLK_FREQ                            ( USER_CLK_FREQ ),
    .USE_RID_PINS                             ( USE_RID_PINS ),
    .VC0_CPL_INFINITE                         ( VC0_CPL_INFINITE ),
    .VC0_RX_RAM_LIMIT                         ( VC0_RX_RAM_LIMIT ),
    .VC0_TOTAL_CREDITS_CD                     ( VC0_TOTAL_CREDITS_CD ),
    .VC0_TOTAL_CREDITS_CH                     ( VC0_TOTAL_CREDITS_CH ),
    .VC0_TOTAL_CREDITS_NPD                    ( VC0_TOTAL_CREDITS_NPD),
    .VC0_TOTAL_CREDITS_NPH                    ( VC0_TOTAL_CREDITS_NPH ),
    .VC0_TOTAL_CREDITS_PD                     ( VC0_TOTAL_CREDITS_PD ),
    .VC0_TOTAL_CREDITS_PH                     ( VC0_TOTAL_CREDITS_PH ),
    .VC0_TX_LASTPACKET                        ( VC0_TX_LASTPACKET ),
    .VC_BASE_PTR                              ( VC_BASE_PTR ),
    .VC_CAP_ID                                ( VC_CAP_ID ),
    .VC_CAP_NEXTPTR                           ( VC_CAP_NEXTPTR ),
    .VC_CAP_ON                                ( VC_CAP_ON ),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS         ( VC_CAP_REJECT_SNOOP_TRANSACTIONS ),
    .VC_CAP_VERSION                           ( VC_CAP_VERSION ),
    .VSEC_BASE_PTR                            ( VSEC_BASE_PTR ),
    .VSEC_CAP_HDR_ID                          ( VSEC_CAP_HDR_ID ),
    .VSEC_CAP_HDR_LENGTH                      ( VSEC_CAP_HDR_LENGTH ),
    .VSEC_CAP_HDR_REVISION                    ( VSEC_CAP_HDR_REVISION ),
    .VSEC_CAP_ID                              ( VSEC_CAP_ID ),
    .VSEC_CAP_IS_LINK_VISIBLE                 ( VSEC_CAP_IS_LINK_VISIBLE ),
    .VSEC_CAP_NEXTPTR                         ( VSEC_CAP_NEXTPTR ),
    .VSEC_CAP_ON                              ( VSEC_CAP_ON ),
    .VSEC_CAP_VERSION                         ( VSEC_CAP_VERSION )
    // I/O
  ) model_ap2_tst_pcie_top_i (

    // AXI Interface
    .user_clk_out                               ( user_clk_out ),
    .user_reset                                 ( bridge_reset_d ),
    .user_lnk_up                                ( user_lnk_up ),

    .user_rst_n                                 ( user_rst_n ),
    .trn_lnk_up                                 ( trn_lnk_up ),

    .tx_buf_av                                  ( tx_buf_av ),
    .tx_err_drop                                ( tx_err_drop ),
    .tx_cfg_req                                 ( tx_cfg_req ),
    .s_axis_tx_tready                           ( s_axis_tx_tready ),
    .s_axis_tx_tdata                            ( s_axis_tx_tdata ),
    .s_axis_tx_tkeep                            ( s_axis_tx_tkeep  ),
    .s_axis_tx_tuser                            ( s_axis_tx_tuser ),
    .s_axis_tx_tlast                            ( s_axis_tx_tlast ),
    .s_axis_tx_tvalid                           ( s_axis_tx_tvalid ),
    .tx_cfg_gnt                                 ( tx_cfg_gnt ),

    .m_axis_rx_tdata                            ( m_axis_rx_tdata ),
    .m_axis_rx_tkeep                            ( m_axis_rx_tkeep ),
    .m_axis_rx_tlast                            ( m_axis_rx_tlast ),
    .m_axis_rx_tvalid                           ( m_axis_rx_tvalid ),
    .m_axis_rx_tready                           ( m_axis_rx_tready ),
    .m_axis_rx_tuser                            ( m_axis_rx_tuser ),
    .rx_np_ok                                   ( rx_np_ok ),
    .rx_np_req                                  ( rx_np_req ),

    .fc_cpld                                    ( fc_cpld ),
    .fc_cplh                                    ( fc_cplh ),
    .fc_npd                                     ( fc_npd ),
    .fc_nph                                     ( fc_nph ),
    .fc_pd                                      ( fc_pd ),
    .fc_ph                                      ( fc_ph ),
    .fc_sel                                     ( fc_sel ),
    .cfg_turnoff_ok                             ( cfg_turnoff_ok ),
    .cfg_received_func_lvl_rst                  ( cfg_received_func_lvl_rst ),

    .cm_rst_n                                   ( 1'b1 ),
    .func_lvl_rst_n                             ( 1'b1 ),
    .lnk_clk_en                                 ( ),
    .cfg_dev_id                                 ( cfg_dev_id ),
    .cfg_vend_id                                ( cfg_vend_id ),
    .cfg_rev_id                                 ( cfg_rev_id ),
    .cfg_subsys_id                              ( cfg_subsys_id ),
    .cfg_subsys_vend_id                         ( cfg_subsys_vend_id ),
    .cfg_pciecap_interrupt_msgnum               ( cfg_pciecap_interrupt_msgnum ),

    .cfg_bridge_serr_en                         ( cfg_bridge_serr_en ),

    .cfg_command_bus_master_enable              ( ),
    .cfg_command_interrupt_disable              ( ),
    .cfg_command_io_enable                      ( ),
    .cfg_command_mem_enable                     ( ),
    .cfg_command_serr_en                        ( ),
    .cfg_dev_control_aux_power_en               ( ),
    .cfg_dev_control_corr_err_reporting_en      ( ),
    .cfg_dev_control_enable_ro                  ( ),
    .cfg_dev_control_ext_tag_en                 ( ),
    .cfg_dev_control_fatal_err_reporting_en     ( ),
    .cfg_dev_control_max_payload                ( ),
    .cfg_dev_control_max_read_req               ( ),
    .cfg_dev_control_non_fatal_reporting_en     ( ),
    .cfg_dev_control_no_snoop_en                ( ),
    .cfg_dev_control_phantom_en                 ( ),
    .cfg_dev_control_ur_err_reporting_en        ( ),
    .cfg_dev_control2_cpl_timeout_dis           ( ),
    .cfg_dev_control2_cpl_timeout_val           ( ),
    .cfg_dev_control2_ari_forward_en            ( ),
    .cfg_dev_control2_atomic_requester_en       ( ),
    .cfg_dev_control2_atomic_egress_block       ( ),
    .cfg_dev_control2_ido_req_en                ( ),
    .cfg_dev_control2_ido_cpl_en                ( ),
    .cfg_dev_control2_ltr_en                    ( ),
    .cfg_dev_control2_tlp_prefix_block          ( ),
    .cfg_dev_status_corr_err_detected           ( ),
    .cfg_dev_status_fatal_err_detected          ( ),
    .cfg_dev_status_non_fatal_err_detected      ( ),
    .cfg_dev_status_ur_detected                 ( ),

    .cfg_mgmt_do                                ( cfg_mgmt_do ),
    .cfg_err_aer_headerlog_set                  ( cfg_err_aer_headerlog_set ),
    .cfg_err_aer_headerlog                      ( cfg_err_aer_headerlog ),
    .cfg_err_cpl_rdy                            ( cfg_err_cpl_rdy ),
    .cfg_interrupt_do                           ( cfg_interrupt_do ),
    .cfg_interrupt_mmenable                     ( cfg_interrupt_mmenable ),
    .cfg_interrupt_msienable                    ( cfg_interrupt_msienable ),
    .cfg_interrupt_msixenable                   ( cfg_interrupt_msixenable ),
    .cfg_interrupt_msixfm                       ( cfg_interrupt_msixfm ),
    .cfg_interrupt_rdy                          ( cfg_interrupt_rdy ),
    .cfg_link_control_rcb                       ( ),
    .cfg_link_control_aspm_control              ( ),
    .cfg_link_control_auto_bandwidth_int_en     ( ),
    .cfg_link_control_bandwidth_int_en          ( ),
    .cfg_link_control_clock_pm_en               ( ),
    .cfg_link_control_common_clock              ( ),
    .cfg_link_control_extended_sync             ( ),
    .cfg_link_control_hw_auto_width_dis         ( ),
    .cfg_link_control_link_disable              ( ),
    .cfg_link_control_retrain_link              ( ),
    .cfg_link_status_auto_bandwidth_status      ( ),
    .cfg_link_status_bandwidth_status           ( ),
    .cfg_link_status_current_speed              ( ),
    .cfg_link_status_dll_active                 ( ),
    .cfg_link_status_link_training              ( ),
    .cfg_link_status_negotiated_width           ( ),
    .cfg_msg_data                               ( cfg_msg_data ),
    .cfg_msg_received                           ( cfg_msg_received ),
    .cfg_msg_received_assert_int_a              ( cfg_msg_received_assert_int_a ),
    .cfg_msg_received_assert_int_b              ( cfg_msg_received_assert_int_b ),
    .cfg_msg_received_assert_int_c              ( cfg_msg_received_assert_int_c ),
    .cfg_msg_received_assert_int_d              ( cfg_msg_received_assert_int_d ),
    .cfg_msg_received_deassert_int_a            ( cfg_msg_received_deassert_int_a ),
    .cfg_msg_received_deassert_int_b            ( cfg_msg_received_deassert_int_b ),
    .cfg_msg_received_deassert_int_c            ( cfg_msg_received_deassert_int_c ),
    .cfg_msg_received_deassert_int_d            ( cfg_msg_received_deassert_int_d ),
    .cfg_msg_received_err_cor                   ( cfg_msg_received_err_cor ),
    .cfg_msg_received_err_fatal                 ( cfg_msg_received_err_fatal ),
    .cfg_msg_received_err_non_fatal             ( cfg_msg_received_err_non_fatal ),
    .cfg_msg_received_pm_as_nak                 ( cfg_msg_received_pm_as_nak ),
    .cfg_msg_received_pme_to                    ( ),
    .cfg_msg_received_pme_to_ack                ( cfg_msg_received_pme_to_ack ),
    .cfg_msg_received_pm_pme                    ( cfg_msg_received_pm_pme ),
    .cfg_msg_received_setslotpowerlimit         ( cfg_msg_received_setslotpowerlimit ),
    .cfg_msg_received_unlock                    ( ),
    .cfg_to_turnoff                             ( cfg_to_turnoff ),
    .cfg_status                                 ( cfg_status ),
    .cfg_command                                ( cfg_command ),
    .cfg_dstatus                                ( cfg_dstatus ),
    .cfg_dcommand                               ( cfg_dcommand ),
    .cfg_lstatus                                ( cfg_lstatus ),
    .cfg_lcommand                               ( cfg_lcommand ),
    .cfg_dcommand2                              ( cfg_dcommand2 ),
    .cfg_pcie_link_state                        ( cfg_pcie_link_state ),
    .cfg_pmcsr_pme_en                           ( cfg_pmcsr_pme_en ),
    .cfg_pmcsr_powerstate                       ( cfg_pmcsr_powerstate ),
    .cfg_pmcsr_pme_status                       ( cfg_pmcsr_pme_status ),
    .cfg_pm_rcv_as_req_l1_n                     ( ),
    .cfg_pm_rcv_enter_l1_n                      ( ),
    .cfg_pm_rcv_enter_l23_n                     ( ),
    .cfg_pm_rcv_req_ack_n                       ( ),
    .cfg_mgmt_rd_wr_done                        ( cfg_mgmt_rd_wr_done ),
    .cfg_slot_control_electromech_il_ctl_pulse  ( cfg_slot_control_electromech_il_ctl_pulse ),
    .cfg_root_control_syserr_corr_err_en        ( cfg_root_control_syserr_corr_err_en ),
    .cfg_root_control_syserr_non_fatal_err_en   ( cfg_root_control_syserr_non_fatal_err_en ),
    .cfg_root_control_syserr_fatal_err_en       ( cfg_root_control_syserr_fatal_err_en ),
    .cfg_root_control_pme_int_en                ( cfg_root_control_pme_int_en),
    .cfg_aer_ecrc_check_en                      ( cfg_aer_ecrc_check_en ),
    .cfg_aer_ecrc_gen_en                        ( cfg_aer_ecrc_gen_en ),
    .cfg_aer_rooterr_corr_err_reporting_en      ( cfg_aer_rooterr_corr_err_reporting_en ),
    .cfg_aer_rooterr_non_fatal_err_reporting_en ( cfg_aer_rooterr_non_fatal_err_reporting_en ),
    .cfg_aer_rooterr_fatal_err_reporting_en     ( cfg_aer_rooterr_fatal_err_reporting_en ),
    .cfg_aer_rooterr_corr_err_received          ( cfg_aer_rooterr_corr_err_received ),
    .cfg_aer_rooterr_non_fatal_err_received     ( cfg_aer_rooterr_non_fatal_err_received ),
    .cfg_aer_rooterr_fatal_err_received         ( cfg_aer_rooterr_fatal_err_received ),
    .cfg_aer_interrupt_msgnum                   ( cfg_aer_interrupt_msgnum ),
    .cfg_transaction                            ( ),
    .cfg_transaction_addr                       ( ),
    .cfg_transaction_type                       ( ),
    .cfg_vc_tcvc_map                            ( cfg_vc_tcvc_map ),
    .cfg_mgmt_byte_en_n                         ( ~cfg_mgmt_byte_en ),
    .cfg_mgmt_di                                ( cfg_mgmt_di ),
    .cfg_dsn                                    ( cfg_dsn ),
    .cfg_mgmt_dwaddr                            ( cfg_mgmt_dwaddr ),
    .cfg_err_acs_n                              ( 1'b1 ),
    .cfg_err_cor_n                              ( ~cfg_err_cor ),
    .cfg_err_cpl_abort_n                        ( ~cfg_err_cpl_abort ),
    .cfg_err_cpl_timeout_n                      ( ~cfg_err_cpl_timeout ),
    .cfg_err_cpl_unexpect_n                     ( ~cfg_err_cpl_unexpect ),
    .cfg_err_ecrc_n                             ( ~cfg_err_ecrc ),
    .cfg_err_locked_n                           ( ~cfg_err_locked ),
    .cfg_err_posted_n                           ( ~cfg_err_posted ),
    .cfg_err_tlp_cpl_header                     ( cfg_err_tlp_cpl_header ),
    .cfg_err_ur_n                               ( ~cfg_err_ur ),
    .cfg_err_malformed_n                        ( ~cfg_err_malformed ),
    .cfg_err_poisoned_n                         ( ~cfg_err_poisoned ),
    .cfg_err_atomic_egress_blocked_n            ( ~cfg_err_atomic_egress_blocked ),
    .cfg_err_mc_blocked_n                       ( ~cfg_err_mc_blocked ),
    .cfg_err_internal_uncor_n                   ( ~cfg_err_internal_uncor ),
    .cfg_err_internal_cor_n                     ( ~cfg_err_internal_cor ),
    .cfg_err_norecovery_n                       ( ~cfg_err_norecovery ),

    .cfg_interrupt_assert_n                     ( ~cfg_interrupt_assert ),
    .cfg_interrupt_di                           ( cfg_interrupt_di ),
    .cfg_interrupt_n                            ( ~cfg_interrupt ),
    .cfg_interrupt_stat_n                       ( ~cfg_interrupt_stat ),
    .cfg_bus_number                             ( cfg_bus_number ),
    .cfg_device_number                          ( cfg_device_number ),
    .cfg_function_number                        ( cfg_function_number ),
    .cfg_ds_bus_number                          ( cfg_ds_bus_number ),
    .cfg_ds_device_number                       ( cfg_ds_device_number ),
    .cfg_ds_function_number                     ( cfg_ds_function_number ),
    .cfg_pm_send_pme_to_n                       ( 1'b1 ),
    .cfg_pm_wake_n                              ( ~cfg_pm_wake ),
    .cfg_pm_halt_aspm_l0s_n                     ( ~cfg_pm_halt_aspm_l0s ),
    .cfg_pm_halt_aspm_l1_n                      ( ~cfg_pm_halt_aspm_l1 ),
    .cfg_pm_force_state_en_n                    ( ~cfg_pm_force_state_en),
    .cfg_pm_force_state                         ( cfg_pm_force_state ),
    .cfg_force_mps                              ( 3'b0 ),
    .cfg_force_common_clock_off                 ( 1'b0 ),
    .cfg_force_extended_sync_on                 ( 1'b0 ),
    .cfg_port_number                            ( 8'b0 ),
    .cfg_mgmt_rd_en_n                           ( ~cfg_mgmt_rd_en ),
    .cfg_trn_pending                            ( cfg_trn_pending ),
    .cfg_mgmt_wr_en_n                           ( ~cfg_mgmt_wr_en ),
    .cfg_mgmt_wr_readonly_n                     ( ~cfg_mgmt_wr_readonly ),
    .cfg_mgmt_wr_rw1c_as_rw_n                   ( ~cfg_mgmt_wr_rw1c_as_rw ),

    .pl_initial_link_width                      ( pl_initial_link_width ),
    .pl_lane_reversal_mode                      ( pl_lane_reversal_mode ),
    .pl_link_gen2_cap                           ( pl_link_gen2_cap ),
    .pl_link_partner_gen2_supported             ( pl_link_partner_gen2_supported ),
    .pl_link_upcfg_cap                          ( pl_link_upcfg_cap ),
    .pl_ltssm_state                             ( pl_ltssm_state_int ),
    .pl_phy_lnk_up                              ( pl_phy_lnk_up_wire ),
    .pl_received_hot_rst                        ( pl_received_hot_rst_wire ),
    .pl_rx_pm_state                             ( pl_rx_pm_state ),
    .pl_sel_lnk_rate                            ( pl_sel_lnk_rate ),
    .pl_sel_lnk_width                           ( pl_sel_lnk_width ),
    .pl_tx_pm_state                             ( pl_tx_pm_state ),
    .pl_directed_link_auton                     ( pl_directed_link_auton ),
    .pl_directed_link_change                    ( pl_directed_link_change ),
    .pl_directed_link_speed                     ( pl_directed_link_speed ),
    .pl_directed_link_width                     ( pl_directed_link_width ),
    .pl_downstream_deemph_source                ( pl_downstream_deemph_source ),
    .pl_upstream_prefer_deemph                  ( pl_upstream_prefer_deemph ),
    .pl_transmit_hot_rst                        ( pl_transmit_hot_rst ),
    .pl_directed_ltssm_new_vld                  ( 1'b0 ),
    .pl_directed_ltssm_new                      ( 6'b0 ),
    .pl_directed_ltssm_stall                    ( 1'b0 ),
    .pl_directed_change_done                    ( pl_directed_change_done ),

    .phy_rdy_n                                  ( phy_rdy_n ),
    .dbg_sclr_a                                 ( ),
    .dbg_sclr_b                                 ( ),
    .dbg_sclr_c                                 ( ),
    .dbg_sclr_d                                 ( ),
    .dbg_sclr_e                                 ( ),
    .dbg_sclr_f                                 ( ),
    .dbg_sclr_g                                 ( ),
    .dbg_sclr_h                                 ( ),
    .dbg_sclr_i                                 ( ),
    .dbg_sclr_j                                 ( ),
    .dbg_sclr_k                                 ( ),

    .dbg_vec_a                                  ( ),
    .dbg_vec_b                                  ( ),
    .dbg_vec_c                                  ( ),
    .pl_dbg_vec                                 ( ),
    .trn_rdllp_data                             ( ),
    .trn_rdllp_src_rdy                          ( ),
    .dbg_mode                                   ( ),
    .dbg_sub_mode                               ( ),
    .pl_dbg_mode                                ( ),

    .drp_clk                                    ( 1'b0 ),
    .drp_do                                     (  ),
    .drp_rdy                                    (  ),
    .drp_addr                                   ( 9'b0 ),
    .drp_en                                     ( 1'b0 ),
    .drp_di                                     ( 16'b0 ),
    .drp_we                                     ( 1'b0 ),

    // Pipe Interface

    .pipe_clk                                   ( pipe_clk            ),
    .user_clk                                   ( user_clk            ),
    .user_clk2                                  ( user_clk2           ),
    .pipe_rx0_polarity_gt                       ( pipe_rx0_polarity_gt       ),
    .pipe_rx1_polarity_gt                       ( pipe_rx1_polarity_gt       ),
    .pipe_rx2_polarity_gt                       ( pipe_rx2_polarity_gt       ),
    .pipe_rx3_polarity_gt                       ( pipe_rx3_polarity_gt       ),
    .pipe_rx4_polarity_gt                       ( pipe_rx4_polarity_gt       ),
    .pipe_rx5_polarity_gt                       ( pipe_rx5_polarity_gt       ),
    .pipe_rx6_polarity_gt                       ( pipe_rx6_polarity_gt       ),
    .pipe_rx7_polarity_gt                       ( pipe_rx7_polarity_gt       ),
    .pipe_tx_deemph_gt                          ( pipe_tx_deemph_gt          ),
    .pipe_tx_margin_gt                          ( pipe_tx_margin_gt          ),
    .pipe_tx_rate_gt                            ( pipe_tx_rate_gt            ),
    .pipe_tx_rcvr_det_gt                        ( pipe_tx_rcvr_det_gt        ),
    .pipe_tx0_char_is_k_gt                      ( pipe_tx0_char_is_k_gt      ),
    .pipe_tx0_compliance_gt                     ( pipe_tx0_compliance_gt     ),
    .pipe_tx0_data_gt                           ( pipe_tx0_data_gt           ),
    .pipe_tx0_elec_idle_gt                      ( pipe_tx0_elec_idle_gt      ),
    .pipe_tx0_powerdown_gt                      ( pipe_tx0_powerdown_gt      ),
    .pipe_tx1_char_is_k_gt                      ( pipe_tx1_char_is_k_gt      ),
    .pipe_tx1_compliance_gt                     ( pipe_tx1_compliance_gt     ),
    .pipe_tx1_data_gt                           ( pipe_tx1_data_gt           ),
    .pipe_tx1_elec_idle_gt                      ( pipe_tx1_elec_idle_gt      ),
    .pipe_tx1_powerdown_gt                      ( pipe_tx1_powerdown_gt      ),
    .pipe_tx2_char_is_k_gt                      ( pipe_tx2_char_is_k_gt      ),
    .pipe_tx2_compliance_gt                     ( pipe_tx2_compliance_gt     ),
    .pipe_tx2_data_gt                           ( pipe_tx2_data_gt           ),
    .pipe_tx2_elec_idle_gt                      ( pipe_tx2_elec_idle_gt      ),
    .pipe_tx2_powerdown_gt                      ( pipe_tx2_powerdown_gt      ),
    .pipe_tx3_char_is_k_gt                      ( pipe_tx3_char_is_k_gt      ),
    .pipe_tx3_compliance_gt                     ( pipe_tx3_compliance_gt     ),
    .pipe_tx3_data_gt                           ( pipe_tx3_data_gt           ),
    .pipe_tx3_elec_idle_gt                      ( pipe_tx3_elec_idle_gt      ),
    .pipe_tx3_powerdown_gt                      ( pipe_tx3_powerdown_gt      ),
    .pipe_tx4_char_is_k_gt                      ( pipe_tx4_char_is_k_gt      ),
    .pipe_tx4_compliance_gt                     ( pipe_tx4_compliance_gt     ),
    .pipe_tx4_data_gt                           ( pipe_tx4_data_gt           ),
    .pipe_tx4_elec_idle_gt                      ( pipe_tx4_elec_idle_gt      ),
    .pipe_tx4_powerdown_gt                      ( pipe_tx4_powerdown_gt      ),
    .pipe_tx5_char_is_k_gt                      ( pipe_tx5_char_is_k_gt      ),
    .pipe_tx5_compliance_gt                     ( pipe_tx5_compliance_gt     ),
    .pipe_tx5_data_gt                           ( pipe_tx5_data_gt           ),
    .pipe_tx5_elec_idle_gt                      ( pipe_tx5_elec_idle_gt      ),
    .pipe_tx5_powerdown_gt                      ( pipe_tx5_powerdown_gt      ),
    .pipe_tx6_char_is_k_gt                      ( pipe_tx6_char_is_k_gt      ),
    .pipe_tx6_compliance_gt                     ( pipe_tx6_compliance_gt     ),
    .pipe_tx6_data_gt                           ( pipe_tx6_data_gt           ),
    .pipe_tx6_elec_idle_gt                      ( pipe_tx6_elec_idle_gt      ),
    .pipe_tx6_powerdown_gt                      ( pipe_tx6_powerdown_gt      ),
    .pipe_tx7_char_is_k_gt                      ( pipe_tx7_char_is_k_gt      ),
    .pipe_tx7_compliance_gt                     ( pipe_tx7_compliance_gt     ),
    .pipe_tx7_data_gt                           ( pipe_tx7_data_gt           ),
    .pipe_tx7_elec_idle_gt                      ( pipe_tx7_elec_idle_gt      ),
    .pipe_tx7_powerdown_gt                      ( pipe_tx7_powerdown_gt      ),

    .pipe_rx0_chanisaligned_gt                  ( pipe_rx0_chanisaligned_gt  ),
    .pipe_rx0_char_is_k_gt                      ( pipe_rx0_char_is_k_gt      ),
    .pipe_rx0_data_gt                           ( pipe_rx0_data_gt           ),
    .pipe_rx0_elec_idle_gt                      ( pipe_rx0_elec_idle_gt      ),
    .pipe_rx0_phy_status_gt                     ( pipe_rx0_phy_status_gt     ),
    .pipe_rx0_status_gt                         ( pipe_rx0_status_gt         ),
    .pipe_rx0_valid_gt                          ( pipe_rx0_valid_gt          ),
    .pipe_rx1_chanisaligned_gt                  ( pipe_rx1_chanisaligned_gt  ),
    .pipe_rx1_char_is_k_gt                      ( pipe_rx1_char_is_k_gt      ),
    .pipe_rx1_data_gt                           ( pipe_rx1_data_gt           ),
    .pipe_rx1_elec_idle_gt                      ( pipe_rx1_elec_idle_gt      ),
    .pipe_rx1_phy_status_gt                     ( pipe_rx1_phy_status_gt     ),
    .pipe_rx1_status_gt                         ( pipe_rx1_status_gt         ),
    .pipe_rx1_valid_gt                          ( pipe_rx1_valid_gt          ),
    .pipe_rx2_chanisaligned_gt                  ( pipe_rx2_chanisaligned_gt  ),
    .pipe_rx2_char_is_k_gt                      ( pipe_rx2_char_is_k_gt      ),
    .pipe_rx2_data_gt                           ( pipe_rx2_data_gt           ),
    .pipe_rx2_elec_idle_gt                      ( pipe_rx2_elec_idle_gt      ),
    .pipe_rx2_phy_status_gt                     ( pipe_rx2_phy_status_gt     ),
    .pipe_rx2_status_gt                         ( pipe_rx2_status_gt         ),
    .pipe_rx2_valid_gt                          ( pipe_rx2_valid_gt          ),
    .pipe_rx3_chanisaligned_gt                  ( pipe_rx3_chanisaligned_gt  ),
    .pipe_rx3_char_is_k_gt                      ( pipe_rx3_char_is_k_gt      ),
    .pipe_rx3_data_gt                           ( pipe_rx3_data_gt           ),
    .pipe_rx3_elec_idle_gt                      ( pipe_rx3_elec_idle_gt      ),
    .pipe_rx3_phy_status_gt                     ( pipe_rx3_phy_status_gt     ),
    .pipe_rx3_status_gt                         ( pipe_rx3_status_gt         ),
    .pipe_rx3_valid_gt                          ( pipe_rx3_valid_gt          ),
    .pipe_rx4_chanisaligned_gt                  ( pipe_rx4_chanisaligned_gt  ),
    .pipe_rx4_char_is_k_gt                      ( pipe_rx4_char_is_k_gt      ),
    .pipe_rx4_data_gt                           ( pipe_rx4_data_gt           ),
    .pipe_rx4_elec_idle_gt                      ( pipe_rx4_elec_idle_gt      ),
    .pipe_rx4_phy_status_gt                     ( pipe_rx4_phy_status_gt     ),
    .pipe_rx4_status_gt                         ( pipe_rx4_status_gt         ),
    .pipe_rx4_valid_gt                          ( pipe_rx4_valid_gt          ),
    .pipe_rx5_chanisaligned_gt                  ( pipe_rx5_chanisaligned_gt  ),
    .pipe_rx5_char_is_k_gt                      ( pipe_rx5_char_is_k_gt      ),
    .pipe_rx5_data_gt                           ( pipe_rx5_data_gt           ),
    .pipe_rx5_elec_idle_gt                      ( pipe_rx5_elec_idle_gt      ),
    .pipe_rx5_phy_status_gt                     ( pipe_rx5_phy_status_gt     ),
    .pipe_rx5_status_gt                         ( pipe_rx5_status_gt         ),
    .pipe_rx5_valid_gt                          ( pipe_rx5_valid_gt          ),
    .pipe_rx6_chanisaligned_gt                  ( pipe_rx6_chanisaligned_gt  ),
    .pipe_rx6_char_is_k_gt                      ( pipe_rx6_char_is_k_gt      ),
    .pipe_rx6_data_gt                           ( pipe_rx6_data_gt           ),
    .pipe_rx6_elec_idle_gt                      ( pipe_rx6_elec_idle_gt      ),
    .pipe_rx6_phy_status_gt                     ( pipe_rx6_phy_status_gt     ),
    .pipe_rx6_status_gt                         ( pipe_rx6_status_gt         ),
    .pipe_rx6_valid_gt                          ( pipe_rx6_valid_gt          ),
    .pipe_rx7_chanisaligned_gt                  ( pipe_rx7_chanisaligned_gt  ),
    .pipe_rx7_char_is_k_gt                      ( pipe_rx7_char_is_k_gt      ),
    .pipe_rx7_data_gt                           ( pipe_rx7_data_gt           ),
    .pipe_rx7_elec_idle_gt                      ( pipe_rx7_elec_idle_gt      ),
    .pipe_rx7_phy_status_gt                     ( pipe_rx7_phy_status_gt     ),
    .pipe_rx7_status_gt                         ( pipe_rx7_status_gt         ),
    .pipe_rx7_valid_gt                          ( pipe_rx7_valid_gt          )

  );
  assign  common_commands_out = 12'b0;  
  assign  pipe_tx_0_sigs      = 25'b0;   
  assign  pipe_tx_1_sigs      = 25'b0; 
  assign  pipe_tx_2_sigs      = 25'b0; 
  assign  pipe_tx_3_sigs      = 25'b0; 
  assign  pipe_tx_4_sigs      = 25'b0; 
  assign  pipe_tx_5_sigs      = 25'b0; 
  assign  pipe_tx_6_sigs      = 25'b0; 
  assign  pipe_tx_7_sigs      = 25'b0; 
end
else
begin
  //------------------------------------------------------------------------------------------------------------------//
  // **** PCI Express Core Wrapper ****                                                                               //
  // The PCI Express Core Wrapper includes the following:                                                             //
  //   1) AXI Streaming Bridge                                                                                        //
  //   2) PCIE 2_1 Hard Block                                                                                         //
  //   3) PCIE PIPE Interface Pipeline                                                                                //
  //------------------------------------------------------------------------------------------------------------------//
  
  /////////////// phy_rdy, rcvr det , speed_change & gt_powerdown /////////////////////////////
    localparam USERCLK2_FREQ     = (USER_CLK2_DIV2 == "TRUE") ? (USER_CLK_FREQ == 4) ? 3 : (USER_CLK_FREQ == 3) ? 2 : USER_CLK_FREQ: USER_CLK_FREQ;
   
    reg [31:0] phy_rdy_reg = 32'b0;
    reg [31:0] rcvr_det_reg     = 32'b0;
    reg  [2:0] pipe_rate_reg    = 3'b0;
    reg  [7:0] gt_powerdown_reg = {4{2'b10}};
    
    wire      rcvr_det;
    wire      speed_change;
    wire      gt_powerdown;
    wire      phy_rdy;
      
    always @ (posedge pipe_clk)
    begin
     phy_rdy_reg      <= {phy_rdy_reg[30:0], sys_rst_n};
     rcvr_det_reg     <= {rcvr_det_reg[30:0], pipe_tx_rcvr_det_gt};
     pipe_rate_reg    <= {pipe_rate_reg[2:0], common_commands_out[1]};
     gt_powerdown_reg <= {gt_powerdown_reg[5:0],pipe_tx_0_sigs[22:21]};
    end 
    
    assign pipe_tx_0_sigs[24:23] = 2'b00;
    assign pipe_tx_1_sigs[24:23] = 2'b00;
    assign pipe_tx_2_sigs[24:23] = 2'b00;
    assign pipe_tx_3_sigs[24:23] = 2'b00;
    assign pipe_tx_4_sigs[24:23] = 2'b00;
    assign pipe_tx_5_sigs[24:23] = 2'b00;
    assign pipe_tx_6_sigs[24:23] = 2'b00;
    assign pipe_tx_7_sigs[24:23] = 2'b00;
    assign phy_rdy      =  phy_rdy_reg[31];
    assign rcvr_det     =  ~rcvr_det_reg[30] && rcvr_det_reg[29];
    assign speed_change = (pipe_rate_reg[2] != pipe_rate_reg[1])? 1'b1 : 1'b0;
    assign gt_powerdown = (gt_powerdown_reg[7:6] == 2'b10 && gt_powerdown_reg[5:4] == 2'b0)? 1'b1 : 1'b0;
    
    //////// generate Rx status and Phy status ////////////// 
    
    wire [2:0] rx_status;
    wire       phy_status;
    
    assign  rx_status  = (pipe_tx_rcvr_det_gt && rcvr_det) ? 3'b011 : 3'b0;
    assign  phy_status = (pipe_tx_rcvr_det_gt && rcvr_det) || speed_change || gt_powerdown ;
  
    //////// generate clocks for pipe mode //////////////
   
    wire clk_500;
    wire clk_250;
    wire clk_125;
    wire clk_62_5;
   
    sys_clk_gen     #(.offset(7000),.halfcycle(1000)) clk_gen_500  (.sys_clk(clk_500));
    sys_clk_gen     #(.offset(6000),.halfcycle(2000)) clk_gen_250  (.sys_clk(clk_250));
    sys_clk_gen     #(.offset(4000),.halfcycle(4000)) clk_gen_125  (.sys_clk(clk_125));
    sys_clk_gen     #(.offset(0000),.halfcycle(8000)) clk_gen_62_5 (.sys_clk(clk_62_5));
   
  
    assign pipe_clk = common_commands_in[0];
    assign user_clk = (USER_CLK_FREQ == 4) ? clk_500 : (USER_CLK_FREQ == 3) ? clk_250 : (USER_CLK_FREQ == 2) ? clk_125 : clk_62_5;
    assign user_clk2 = (USERCLK2_FREQ == 4) ? clk_500 : (USERCLK2_FREQ == 3) ? clk_250 : (USERCLK2_FREQ == 2) ? clk_125 : clk_62_5;
    
model_ap2_tst_pcie_top # (
    .PIPE_PIPELINE_STAGES                     ( PIPE_PIPELINE_STAGES ),
    .AER_BASE_PTR                             ( AER_BASE_PTR ),
    .AER_CAP_ECRC_CHECK_CAPABLE               ( AER_CAP_ECRC_CHECK_CAPABLE ),
    .AER_CAP_ECRC_GEN_CAPABLE                 ( AER_CAP_ECRC_GEN_CAPABLE ),
    .AER_CAP_ID                               ( AER_CAP_ID ),
    .AER_CAP_MULTIHEADER                      ( AER_CAP_MULTIHEADER ),
    .AER_CAP_NEXTPTR                          ( AER_CAP_NEXTPTR ),
    .AER_CAP_ON                               ( AER_CAP_ON ),
    .AER_CAP_OPTIONAL_ERR_SUPPORT             ( AER_CAP_OPTIONAL_ERR_SUPPORT ),
    .AER_CAP_PERMIT_ROOTERR_UPDATE            ( AER_CAP_PERMIT_ROOTERR_UPDATE ),
    .AER_CAP_VERSION                          ( AER_CAP_VERSION ),
    .ALLOW_X8_GEN2                            ( ALLOW_X8_GEN2 ),
    .BAR0                                     ( BAR0 ),
    .BAR1                                     ( BAR1 ),
    .BAR2                                     ( BAR2 ),
    .BAR3                                     ( BAR3 ),
    .BAR4                                     ( BAR4 ),
    .BAR5                                     ( BAR5 ),
    .C_DATA_WIDTH                             ( C_DATA_WIDTH ),
    .CAPABILITIES_PTR                         ( CAPABILITIES_PTR ),
    .CARDBUS_CIS_POINTER                      ( CARDBUS_CIS_POINTER ),
    .CFG_ECRC_ERR_CPLSTAT                     ( CFG_ECRC_ERR_CPLSTAT ),
    .CLASS_CODE                               ( CLASS_CODE ),
    .CMD_INTX_IMPLEMENTED                     ( CMD_INTX_IMPLEMENTED ),
    .CPL_TIMEOUT_DISABLE_SUPPORTED            ( CPL_TIMEOUT_DISABLE_SUPPORTED ),
    .CPL_TIMEOUT_RANGES_SUPPORTED             ( CPL_TIMEOUT_RANGES_SUPPORTED ),
    .CRM_MODULE_RSTS                          ( CRM_MODULE_RSTS ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE ),
    .DEV_CAP_ENDPOINT_L0S_LATENCY             ( DEV_CAP_ENDPOINT_L0S_LATENCY ),
    .DEV_CAP_ENDPOINT_L1_LATENCY              ( DEV_CAP_ENDPOINT_L1_LATENCY ),
    .DEV_CAP_EXT_TAG_SUPPORTED                ( DEV_CAP_EXT_TAG_SUPPORTED ),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     ( DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE ),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED            ( DEV_CAP_MAX_PAYLOAD_SUPPORTED ),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        ( DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT ),
    .DEV_CAP_ROLE_BASED_ERROR                 ( DEV_CAP_ROLE_BASED_ERROR ),
    .DEV_CAP_RSVD_14_12                       ( DEV_CAP_RSVD_14_12 ),
    .DEV_CAP_RSVD_17_16                       ( DEV_CAP_RSVD_17_16 ),
    .DEV_CAP_RSVD_31_29                       ( DEV_CAP_RSVD_31_29 ),
    .DEV_CONTROL_AUX_POWER_SUPPORTED          ( DEV_CONTROL_AUX_POWER_SUPPORTED ),
    .DEV_CONTROL_EXT_TAG_DEFAULT              ( DEV_CONTROL_EXT_TAG_DEFAULT ),
    .DISABLE_ASPM_L1_TIMER                    ( DISABLE_ASPM_L1_TIMER ),
    .DISABLE_BAR_FILTERING                    ( DISABLE_BAR_FILTERING ),
    .DISABLE_ID_CHECK                         ( DISABLE_ID_CHECK ),
    .DISABLE_LANE_REVERSAL                    ( DISABLE_LANE_REVERSAL ),
    .DISABLE_RX_POISONED_RESP                 ( DISABLE_RX_POISONED_RESP ),
    .DISABLE_RX_TC_FILTER                     ( DISABLE_RX_TC_FILTER ),
    .DISABLE_SCRAMBLING                       ( DISABLE_SCRAMBLING ),
    .DNSTREAM_LINK_NUM                        ( DNSTREAM_LINK_NUM ),
    .DSN_BASE_PTR                             ( DSN_BASE_PTR ),
    .DSN_CAP_ID                               ( DSN_CAP_ID ),
    .DSN_CAP_NEXTPTR                          ( DSN_CAP_NEXTPTR ),
    .DSN_CAP_ON                               ( DSN_CAP_ON ),
    .DSN_CAP_VERSION                          ( DSN_CAP_VERSION ),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED        ( DEV_CAP2_ARI_FORWARDING_SUPPORTED ),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      ( DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED ),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED      ( DEV_CAP2_CAS128_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     ( DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED ),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    ( DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED ),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED         ( DEV_CAP2_LTR_MECHANISM_SUPPORTED ),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         ( DEV_CAP2_MAX_ENDEND_TLP_PREFIXES ),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      ( DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING ),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED         ( DEV_CAP2_TPH_COMPLETER_SUPPORTED ),
    .DISABLE_ERR_MSG                          ( DISABLE_ERR_MSG ),
    .DISABLE_LOCKED_FILTER                    ( DISABLE_LOCKED_FILTER ),
    .DISABLE_PPM_FILTER                       ( DISABLE_PPM_FILTER ),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   ( ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED ),
    .ENABLE_MSG_ROUTE                         ( ENABLE_MSG_ROUTE ),
    .ENABLE_RX_TD_ECRC_TRIM                   ( ENABLE_RX_TD_ECRC_TRIM ),
    .ENTER_RVRY_EI_L0                         ( ENTER_RVRY_EI_L0 ),
    .EXIT_LOOPBACK_ON_EI                      ( EXIT_LOOPBACK_ON_EI ),
    .EXPANSION_ROM                            ( EXPANSION_ROM ),
    .EXT_CFG_CAP_PTR                          ( EXT_CFG_CAP_PTR ),
    .EXT_CFG_XP_CAP_PTR                       ( EXT_CFG_XP_CAP_PTR ),
    .HEADER_TYPE                              ( HEADER_TYPE ),
    .INFER_EI                                 ( INFER_EI ),
    .INTERRUPT_PIN                            ( INTERRUPT_PIN ),
    .INTERRUPT_STAT_AUTO                      ( INTERRUPT_STAT_AUTO ),
    .IS_SWITCH                                ( IS_SWITCH ),
    .LAST_CONFIG_DWORD                        ( LAST_CONFIG_DWORD ),
    .LINK_CAP_ASPM_OPTIONALITY                ( LINK_CAP_ASPM_OPTIONALITY ),
    .LINK_CAP_ASPM_SUPPORT                    ( LINK_CAP_ASPM_SUPPORT ),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT          ( LINK_CAP_CLOCK_POWER_MANAGEMENT ),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   ( LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1           ( LINK_CAP_L0S_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2           ( LINK_CAP_L0S_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1            ( LINK_CAP_L1_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2            ( LINK_CAP_L1_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ( LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ),
    .LINK_CAP_MAX_LINK_SPEED                  ( LINK_CAP_MAX_LINK_SPEED ),
    .LINK_CAP_MAX_LINK_WIDTH                  ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_RSVD_23                         ( LINK_CAP_RSVD_23 ),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     ( LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE ),
    .LINK_CONTROL_RCB                         ( LINK_CONTROL_RCB ),
    .LINK_CTRL2_DEEMPHASIS                    ( LINK_CTRL2_DEEMPHASIS ),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   ( LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE ),
    .LINK_CTRL2_TARGET_LINK_SPEED             ( LINK_CTRL2_TARGET_LINK_SPEED ),
    .LINK_STATUS_SLOT_CLOCK_CONFIG            ( LINK_STATUS_SLOT_CLOCK_CONFIG ),
    .LL_ACK_TIMEOUT                           ( LL_ACK_TIMEOUT ),
    .LL_ACK_TIMEOUT_EN                        ( LL_ACK_TIMEOUT_EN ),
    .LL_ACK_TIMEOUT_FUNC                      ( LL_ACK_TIMEOUT_FUNC ),
    .LL_REPLAY_TIMEOUT                        ( LL_REPLAY_TIMEOUT ),
    .LL_REPLAY_TIMEOUT_EN                     ( LL_REPLAY_TIMEOUT_EN ),
    .LL_REPLAY_TIMEOUT_FUNC                   ( LL_REPLAY_TIMEOUT_FUNC ),
    .LTSSM_MAX_LINK_WIDTH                     ( LTSSM_MAX_LINK_WIDTH ),
    .MPS_FORCE                                ( MPS_FORCE),
    .MSI_BASE_PTR                             ( MSI_BASE_PTR ),
    .MSI_CAP_ID                               ( MSI_CAP_ID ),
    .MSI_CAP_MULTIMSGCAP                      ( MSI_CAP_MULTIMSGCAP ),
    .MSI_CAP_MULTIMSG_EXTENSION               ( MSI_CAP_MULTIMSG_EXTENSION ),
    .MSI_CAP_NEXTPTR                          ( MSI_CAP_NEXTPTR ),
    .MSI_CAP_ON                               ( MSI_CAP_ON ),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE       ( MSI_CAP_PER_VECTOR_MASKING_CAPABLE ),
    .MSI_CAP_64_BIT_ADDR_CAPABLE              ( MSI_CAP_64_BIT_ADDR_CAPABLE ),
    .MSIX_BASE_PTR                            ( MSIX_BASE_PTR ),
    .MSIX_CAP_ID                              ( MSIX_CAP_ID ),
    .MSIX_CAP_NEXTPTR                         ( MSIX_CAP_NEXTPTR ),
    .MSIX_CAP_ON                              ( MSIX_CAP_ON ),
    .MSIX_CAP_PBA_BIR                         ( MSIX_CAP_PBA_BIR ),
    .MSIX_CAP_PBA_OFFSET                      ( MSIX_CAP_PBA_OFFSET ),
    .MSIX_CAP_TABLE_BIR                       ( MSIX_CAP_TABLE_BIR ),
    .MSIX_CAP_TABLE_OFFSET                    ( MSIX_CAP_TABLE_OFFSET ),
    .MSIX_CAP_TABLE_SIZE                      ( MSIX_CAP_TABLE_SIZE ),
    .N_FTS_COMCLK_GEN1                        ( N_FTS_COMCLK_GEN1 ),
    .N_FTS_COMCLK_GEN2                        ( N_FTS_COMCLK_GEN2 ),
    .N_FTS_GEN1                               ( N_FTS_GEN1 ),
    .N_FTS_GEN2                               ( N_FTS_GEN2 ),
    .PCIE_BASE_PTR                            ( PCIE_BASE_PTR ),
    .PCIE_CAP_CAPABILITY_ID                   ( PCIE_CAP_CAPABILITY_ID ),
    .PCIE_CAP_CAPABILITY_VERSION              ( PCIE_CAP_CAPABILITY_VERSION ),
    .PCIE_CAP_DEVICE_PORT_TYPE                ( PCIE_CAP_DEVICE_PORT_TYPE ),
    .PCIE_CAP_NEXTPTR                         ( PCIE_CAP_NEXTPTR ),
    .PCIE_CAP_ON                              ( PCIE_CAP_ON ),
    .PCIE_CAP_RSVD_15_14                      ( PCIE_CAP_RSVD_15_14 ),
    .PCIE_CAP_SLOT_IMPLEMENTED                ( PCIE_CAP_SLOT_IMPLEMENTED ),
    .PCIE_REVISION                            ( PCIE_REVISION ),
    .PL_AUTO_CONFIG                           ( PL_AUTO_CONFIG ),
    .PL_FAST_TRAIN                            ( PL_FAST_TRAIN ),
    .PM_ASPML0S_TIMEOUT                       ( PM_ASPML0S_TIMEOUT ),
    .PM_ASPML0S_TIMEOUT_EN                    ( PM_ASPML0S_TIMEOUT_EN ),
    .PM_ASPML0S_TIMEOUT_FUNC                  ( PM_ASPML0S_TIMEOUT_FUNC ),
    .PM_ASPM_FASTEXIT                         ( PM_ASPM_FASTEXIT ),
    .PM_BASE_PTR                              ( PM_BASE_PTR ),
    .PM_CAP_AUXCURRENT                        ( PM_CAP_AUXCURRENT ),
    .PM_CAP_D1SUPPORT                         ( PM_CAP_D1SUPPORT ),
    .PM_CAP_D2SUPPORT                         ( PM_CAP_D2SUPPORT ),
    .PM_CAP_DSI                               ( PM_CAP_DSI ),
    .PM_CAP_ID                                ( PM_CAP_ID ),
    .PM_CAP_NEXTPTR                           ( PM_CAP_NEXTPTR ),
    .PM_CAP_ON                                ( PM_CAP_ON ),
    .PM_CAP_PME_CLOCK                         ( PM_CAP_PME_CLOCK ),
    .PM_CAP_PMESUPPORT                        ( PM_CAP_PMESUPPORT ),
    .PM_CAP_RSVD_04                           ( PM_CAP_RSVD_04 ),
    .PM_CAP_VERSION                           ( PM_CAP_VERSION ),
    .PM_CSR_B2B3                              ( PM_CSR_B2B3 ),
    .PM_CSR_BPCCEN                            ( PM_CSR_BPCCEN ),
    .PM_CSR_NOSOFTRST                         ( PM_CSR_NOSOFTRST ),
    .PM_DATA0                                 ( PM_DATA0 ),
    .PM_DATA1                                 ( PM_DATA1 ),
    .PM_DATA2                                 ( PM_DATA2 ),
    .PM_DATA3                                 ( PM_DATA3 ),
    .PM_DATA4                                 ( PM_DATA4 ),
    .PM_DATA5                                 ( PM_DATA5 ),
    .PM_DATA6                                 ( PM_DATA6 ),
    .PM_DATA7                                 ( PM_DATA7 ),
    .PM_DATA_SCALE0                           ( PM_DATA_SCALE0 ),
    .PM_DATA_SCALE1                           ( PM_DATA_SCALE1 ),
    .PM_DATA_SCALE2                           ( PM_DATA_SCALE2 ),
    .PM_DATA_SCALE3                           ( PM_DATA_SCALE3 ),
    .PM_DATA_SCALE4                           ( PM_DATA_SCALE4 ),
    .PM_DATA_SCALE5                           ( PM_DATA_SCALE5 ),
    .PM_DATA_SCALE6                           ( PM_DATA_SCALE6 ),
    .PM_DATA_SCALE7                           ( PM_DATA_SCALE7 ),
    .PM_MF                                    ( PM_MF ),
    .RBAR_BASE_PTR                            ( RBAR_BASE_PTR ),
    .RBAR_CAP_CONTROL_ENCODEDBAR0             ( RBAR_CAP_CONTROL_ENCODEDBAR0 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR1             ( RBAR_CAP_CONTROL_ENCODEDBAR1 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR2             ( RBAR_CAP_CONTROL_ENCODEDBAR2 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR3             ( RBAR_CAP_CONTROL_ENCODEDBAR3 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR4             ( RBAR_CAP_CONTROL_ENCODEDBAR4 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR5             ( RBAR_CAP_CONTROL_ENCODEDBAR5 ),
    .RBAR_CAP_ID                              ( RBAR_CAP_ID),
    .RBAR_CAP_INDEX0                          ( RBAR_CAP_INDEX0 ),
    .RBAR_CAP_INDEX1                          ( RBAR_CAP_INDEX1 ),
    .RBAR_CAP_INDEX2                          ( RBAR_CAP_INDEX2 ),
    .RBAR_CAP_INDEX3                          ( RBAR_CAP_INDEX3 ),
    .RBAR_CAP_INDEX4                          ( RBAR_CAP_INDEX4 ),
    .RBAR_CAP_INDEX5                          ( RBAR_CAP_INDEX5 ),
    .RBAR_CAP_NEXTPTR                         ( RBAR_CAP_NEXTPTR ),
    .RBAR_CAP_ON                              ( RBAR_CAP_ON ),
    .RBAR_CAP_SUP0                            ( RBAR_CAP_SUP0 ),
    .RBAR_CAP_SUP1                            ( RBAR_CAP_SUP1 ),
    .RBAR_CAP_SUP2                            ( RBAR_CAP_SUP2 ),
    .RBAR_CAP_SUP3                            ( RBAR_CAP_SUP3 ),
    .RBAR_CAP_SUP4                            ( RBAR_CAP_SUP4 ),
    .RBAR_CAP_SUP5                            ( RBAR_CAP_SUP5 ),
    .RBAR_CAP_VERSION                         ( RBAR_CAP_VERSION ),
    .RBAR_NUM                                 ( RBAR_NUM ),
    .RECRC_CHK                                ( RECRC_CHK ),
    .RECRC_CHK_TRIM                           ( RECRC_CHK_TRIM ),
    .ROOT_CAP_CRS_SW_VISIBILITY               ( ROOT_CAP_CRS_SW_VISIBILITY ),
    .RP_AUTO_SPD                              ( RP_AUTO_SPD ),
    .RP_AUTO_SPD_LOOPCNT                      ( RP_AUTO_SPD_LOOPCNT ),
    .SELECT_DLL_IF                            ( SELECT_DLL_IF ),
    .SLOT_CAP_ATT_BUTTON_PRESENT              ( SLOT_CAP_ATT_BUTTON_PRESENT ),
    .SLOT_CAP_ATT_INDICATOR_PRESENT           ( SLOT_CAP_ATT_INDICATOR_PRESENT ),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT          ( SLOT_CAP_ELEC_INTERLOCK_PRESENT ),
    .SLOT_CAP_HOTPLUG_CAPABLE                 ( SLOT_CAP_HOTPLUG_CAPABLE ),
    .SLOT_CAP_HOTPLUG_SURPRISE                ( SLOT_CAP_HOTPLUG_SURPRISE ),
    .SLOT_CAP_MRL_SENSOR_PRESENT              ( SLOT_CAP_MRL_SENSOR_PRESENT ),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        ( SLOT_CAP_NO_CMD_COMPLETED_SUPPORT ),
    .SLOT_CAP_PHYSICAL_SLOT_NUM               ( SLOT_CAP_PHYSICAL_SLOT_NUM ),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT        ( SLOT_CAP_POWER_CONTROLLER_PRESENT ),
    .SLOT_CAP_POWER_INDICATOR_PRESENT         ( SLOT_CAP_POWER_INDICATOR_PRESENT ),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE          ( SLOT_CAP_SLOT_POWER_LIMIT_SCALE ),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE          ( SLOT_CAP_SLOT_POWER_LIMIT_VALUE ),
    .SPARE_BIT0                               ( SPARE_BIT0 ),
    .SPARE_BIT1                               ( SPARE_BIT1 ),
    .SPARE_BIT2                               ( SPARE_BIT2 ),
    .SPARE_BIT3                               ( SPARE_BIT3 ),
    .SPARE_BIT4                               ( SPARE_BIT4 ),
    .SPARE_BIT5                               ( SPARE_BIT5 ),
    .SPARE_BIT6                               ( SPARE_BIT6 ),
    .SPARE_BIT7                               ( SPARE_BIT7 ),
    .SPARE_BIT8                               ( SPARE_BIT8 ),
    .SPARE_BYTE0                              ( SPARE_BYTE0 ),
    .SPARE_BYTE1                              ( SPARE_BYTE1 ),
    .SPARE_BYTE2                              ( SPARE_BYTE2 ),
    .SPARE_BYTE3                              ( SPARE_BYTE3 ),
    .SPARE_WORD0                              ( SPARE_WORD0 ),
    .SPARE_WORD1                              ( SPARE_WORD1 ),
    .SPARE_WORD2                              ( SPARE_WORD2 ),
    .SPARE_WORD3                              ( SPARE_WORD3 ),
    .SSL_MESSAGE_AUTO                         ( SSL_MESSAGE_AUTO ),
    .TECRC_EP_INV                             ( TECRC_EP_INV ),
    .TL_RBYPASS                               ( TL_RBYPASS ),
    .TL_RX_RAM_RADDR_LATENCY                  ( TL_RX_RAM_RADDR_LATENCY ),
    .TL_RX_RAM_RDATA_LATENCY                  ( TL_RX_RAM_RDATA_LATENCY ),
    .TL_RX_RAM_WRITE_LATENCY                  ( TL_RX_RAM_WRITE_LATENCY ),
    .TL_TFC_DISABLE                           ( TL_TFC_DISABLE ),
    .TL_TX_CHECKS_DISABLE                     ( TL_TX_CHECKS_DISABLE ),
    .TL_TX_RAM_RADDR_LATENCY                  ( TL_TX_RAM_RADDR_LATENCY ),
    .TL_TX_RAM_RDATA_LATENCY                  ( TL_TX_RAM_RDATA_LATENCY ),
    .TL_TX_RAM_WRITE_LATENCY                  ( TL_TX_RAM_WRITE_LATENCY ),
    .TRN_DW                                   ( TRN_DW ),
    .TRN_NP_FC                                ( TRN_NP_FC ),
    .UPCONFIG_CAPABLE                         ( UPCONFIG_CAPABLE ),
    .UPSTREAM_FACING                          ( UPSTREAM_FACING ),
    .UR_ATOMIC                                ( UR_ATOMIC ),
    .UR_CFG1                                  ( UR_CFG1 ),
    .UR_INV_REQ                               ( UR_INV_REQ ),
    .UR_PRS_RESPONSE                          ( UR_PRS_RESPONSE ),
    .USER_CLK2_DIV2                           ( USER_CLK2_DIV2 ),
    .USER_CLK_FREQ                            ( USER_CLK_FREQ ),
    .USE_RID_PINS                             ( USE_RID_PINS ),
    .VC0_CPL_INFINITE                         ( VC0_CPL_INFINITE ),
    .VC0_RX_RAM_LIMIT                         ( VC0_RX_RAM_LIMIT ),
    .VC0_TOTAL_CREDITS_CD                     ( VC0_TOTAL_CREDITS_CD ),
    .VC0_TOTAL_CREDITS_CH                     ( VC0_TOTAL_CREDITS_CH ),
    .VC0_TOTAL_CREDITS_NPD                    ( VC0_TOTAL_CREDITS_NPD),
    .VC0_TOTAL_CREDITS_NPH                    ( VC0_TOTAL_CREDITS_NPH ),
    .VC0_TOTAL_CREDITS_PD                     ( VC0_TOTAL_CREDITS_PD ),
    .VC0_TOTAL_CREDITS_PH                     ( VC0_TOTAL_CREDITS_PH ),
    .VC0_TX_LASTPACKET                        ( VC0_TX_LASTPACKET ),
    .VC_BASE_PTR                              ( VC_BASE_PTR ),
    .VC_CAP_ID                                ( VC_CAP_ID ),
    .VC_CAP_NEXTPTR                           ( VC_CAP_NEXTPTR ),
    .VC_CAP_ON                                ( VC_CAP_ON ),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS         ( VC_CAP_REJECT_SNOOP_TRANSACTIONS ),
    .VC_CAP_VERSION                           ( VC_CAP_VERSION ),
    .VSEC_BASE_PTR                            ( VSEC_BASE_PTR ),
    .VSEC_CAP_HDR_ID                          ( VSEC_CAP_HDR_ID ),
    .VSEC_CAP_HDR_LENGTH                      ( VSEC_CAP_HDR_LENGTH ),
    .VSEC_CAP_HDR_REVISION                    ( VSEC_CAP_HDR_REVISION ),
    .VSEC_CAP_ID                              ( VSEC_CAP_ID ),
    .VSEC_CAP_IS_LINK_VISIBLE                 ( VSEC_CAP_IS_LINK_VISIBLE ),
    .VSEC_CAP_NEXTPTR                         ( VSEC_CAP_NEXTPTR ),
    .VSEC_CAP_ON                              ( VSEC_CAP_ON ),
    .VSEC_CAP_VERSION                         ( VSEC_CAP_VERSION )
    // I/O
  ) model_ap2_tst_pcie_top_i (

    // AXI Interface
    .user_clk_out                               ( user_clk_out ),
    .user_reset                                 ( bridge_reset_d ),
    .user_lnk_up                                ( user_lnk_up ),

    .user_rst_n                                 ( user_rst_n ),
    .trn_lnk_up                                 ( trn_lnk_up ),

    .tx_buf_av                                  ( tx_buf_av ),
    .tx_err_drop                                ( tx_err_drop ),
    .tx_cfg_req                                 ( tx_cfg_req ),
    .s_axis_tx_tready                           ( s_axis_tx_tready ),
    .s_axis_tx_tdata                            ( s_axis_tx_tdata ),
    .s_axis_tx_tkeep                            ( s_axis_tx_tkeep  ),
    .s_axis_tx_tuser                            ( s_axis_tx_tuser ),
    .s_axis_tx_tlast                            ( s_axis_tx_tlast ),
    .s_axis_tx_tvalid                           ( s_axis_tx_tvalid ),
    .tx_cfg_gnt                                 ( tx_cfg_gnt ),

    .m_axis_rx_tdata                            ( m_axis_rx_tdata ),
    .m_axis_rx_tkeep                            ( m_axis_rx_tkeep ),
    .m_axis_rx_tlast                            ( m_axis_rx_tlast ),
    .m_axis_rx_tvalid                           ( m_axis_rx_tvalid ),
    .m_axis_rx_tready                           ( m_axis_rx_tready ),
    .m_axis_rx_tuser                            ( m_axis_rx_tuser ),
    .rx_np_ok                                   ( rx_np_ok ),
    .rx_np_req                                  ( rx_np_req ),

    .fc_cpld                                    ( fc_cpld ),
    .fc_cplh                                    ( fc_cplh ),
    .fc_npd                                     ( fc_npd ),
    .fc_nph                                     ( fc_nph ),
    .fc_pd                                      ( fc_pd ),
    .fc_ph                                      ( fc_ph ),
    .fc_sel                                     ( fc_sel ),
    .cfg_turnoff_ok                             ( cfg_turnoff_ok ),
    .cfg_received_func_lvl_rst                  ( cfg_received_func_lvl_rst ),

    .cm_rst_n                                   ( 1'b1 ),
    .func_lvl_rst_n                             ( 1'b1 ),
    .lnk_clk_en                                 ( ),
    .cfg_dev_id                                 ( cfg_dev_id ),
    .cfg_vend_id                                ( cfg_vend_id ),
    .cfg_rev_id                                 ( cfg_rev_id ),
    .cfg_subsys_id                              ( cfg_subsys_id ),
    .cfg_subsys_vend_id                         ( cfg_subsys_vend_id ),
    .cfg_pciecap_interrupt_msgnum               ( cfg_pciecap_interrupt_msgnum ),

    .cfg_bridge_serr_en                         ( cfg_bridge_serr_en ),

    .cfg_command_bus_master_enable              ( ),
    .cfg_command_interrupt_disable              ( ),
    .cfg_command_io_enable                      ( ),
    .cfg_command_mem_enable                     ( ),
    .cfg_command_serr_en                        ( ),
    .cfg_dev_control_aux_power_en               ( ),
    .cfg_dev_control_corr_err_reporting_en      ( ),
    .cfg_dev_control_enable_ro                  ( ),
    .cfg_dev_control_ext_tag_en                 ( ),
    .cfg_dev_control_fatal_err_reporting_en     ( ),
    .cfg_dev_control_max_payload                ( ),
    .cfg_dev_control_max_read_req               ( ),
    .cfg_dev_control_non_fatal_reporting_en     ( ),
    .cfg_dev_control_no_snoop_en                ( ),
    .cfg_dev_control_phantom_en                 ( ),
    .cfg_dev_control_ur_err_reporting_en        ( ),
    .cfg_dev_control2_cpl_timeout_dis           ( ),
    .cfg_dev_control2_cpl_timeout_val           ( ),
    .cfg_dev_control2_ari_forward_en            ( ),
    .cfg_dev_control2_atomic_requester_en       ( ),
    .cfg_dev_control2_atomic_egress_block       ( ),
    .cfg_dev_control2_ido_req_en                ( ),
    .cfg_dev_control2_ido_cpl_en                ( ),
    .cfg_dev_control2_ltr_en                    ( ),
    .cfg_dev_control2_tlp_prefix_block          ( ),
    .cfg_dev_status_corr_err_detected           ( ),
    .cfg_dev_status_fatal_err_detected          ( ),
    .cfg_dev_status_non_fatal_err_detected      ( ),
    .cfg_dev_status_ur_detected                 ( ),

    .cfg_mgmt_do                                ( cfg_mgmt_do ),
    .cfg_err_aer_headerlog_set                  ( cfg_err_aer_headerlog_set ),
    .cfg_err_aer_headerlog                      ( cfg_err_aer_headerlog ),
    .cfg_err_cpl_rdy                            ( cfg_err_cpl_rdy ),
    .cfg_interrupt_do                           ( cfg_interrupt_do ),
    .cfg_interrupt_mmenable                     ( cfg_interrupt_mmenable ),
    .cfg_interrupt_msienable                    ( cfg_interrupt_msienable ),
    .cfg_interrupt_msixenable                   ( cfg_interrupt_msixenable ),
    .cfg_interrupt_msixfm                       ( cfg_interrupt_msixfm ),
    .cfg_interrupt_rdy                          ( cfg_interrupt_rdy ),
    .cfg_link_control_rcb                       ( ),
    .cfg_link_control_aspm_control              ( ),
    .cfg_link_control_auto_bandwidth_int_en     ( ),
    .cfg_link_control_bandwidth_int_en          ( ),
    .cfg_link_control_clock_pm_en               ( ),
    .cfg_link_control_common_clock              ( ),
    .cfg_link_control_extended_sync             ( ),
    .cfg_link_control_hw_auto_width_dis         ( ),
    .cfg_link_control_link_disable              ( ),
    .cfg_link_control_retrain_link              ( ),
    .cfg_link_status_auto_bandwidth_status      ( ),
    .cfg_link_status_bandwidth_status           ( ),
    .cfg_link_status_current_speed              ( ),
    .cfg_link_status_dll_active                 ( ),
    .cfg_link_status_link_training              ( ),
    .cfg_link_status_negotiated_width           ( ),
    .cfg_msg_data                               ( cfg_msg_data ),
    .cfg_msg_received                           ( cfg_msg_received ),
    .cfg_msg_received_assert_int_a              ( cfg_msg_received_assert_int_a ),
    .cfg_msg_received_assert_int_b              ( cfg_msg_received_assert_int_b ),
    .cfg_msg_received_assert_int_c              ( cfg_msg_received_assert_int_c ),
    .cfg_msg_received_assert_int_d              ( cfg_msg_received_assert_int_d ),
    .cfg_msg_received_deassert_int_a            ( cfg_msg_received_deassert_int_a ),
    .cfg_msg_received_deassert_int_b            ( cfg_msg_received_deassert_int_b ),
    .cfg_msg_received_deassert_int_c            ( cfg_msg_received_deassert_int_c ),
    .cfg_msg_received_deassert_int_d            ( cfg_msg_received_deassert_int_d ),
    .cfg_msg_received_err_cor                   ( cfg_msg_received_err_cor ),
    .cfg_msg_received_err_fatal                 ( cfg_msg_received_err_fatal ),
    .cfg_msg_received_err_non_fatal             ( cfg_msg_received_err_non_fatal ),
    .cfg_msg_received_pm_as_nak                 ( cfg_msg_received_pm_as_nak ),
    .cfg_msg_received_pme_to                    ( ),
    .cfg_msg_received_pme_to_ack                ( cfg_msg_received_pme_to_ack ),
    .cfg_msg_received_pm_pme                    ( cfg_msg_received_pm_pme ),
    .cfg_msg_received_setslotpowerlimit         ( cfg_msg_received_setslotpowerlimit ),
    .cfg_msg_received_unlock                    ( ),
    .cfg_to_turnoff                             ( cfg_to_turnoff ),
    .cfg_status                                 ( cfg_status ),
    .cfg_command                                ( cfg_command ),
    .cfg_dstatus                                ( cfg_dstatus ),
    .cfg_dcommand                               ( cfg_dcommand ),
    .cfg_lstatus                                ( cfg_lstatus ),
    .cfg_lcommand                               ( cfg_lcommand ),
    .cfg_dcommand2                              ( cfg_dcommand2 ),
    .cfg_pcie_link_state                        ( cfg_pcie_link_state ),
    .cfg_pmcsr_pme_en                           ( cfg_pmcsr_pme_en ),
    .cfg_pmcsr_powerstate                       ( cfg_pmcsr_powerstate ),
    .cfg_pmcsr_pme_status                       ( cfg_pmcsr_pme_status ),
    .cfg_pm_rcv_as_req_l1_n                     ( ),
    .cfg_pm_rcv_enter_l1_n                      ( ),
    .cfg_pm_rcv_enter_l23_n                     ( ),
    .cfg_pm_rcv_req_ack_n                       ( ),
    .cfg_mgmt_rd_wr_done                        ( cfg_mgmt_rd_wr_done ),
    .cfg_slot_control_electromech_il_ctl_pulse  ( cfg_slot_control_electromech_il_ctl_pulse ),
    .cfg_root_control_syserr_corr_err_en        ( cfg_root_control_syserr_corr_err_en ),
    .cfg_root_control_syserr_non_fatal_err_en   ( cfg_root_control_syserr_non_fatal_err_en ),
    .cfg_root_control_syserr_fatal_err_en       ( cfg_root_control_syserr_fatal_err_en ),
    .cfg_root_control_pme_int_en                ( cfg_root_control_pme_int_en),
    .cfg_aer_ecrc_check_en                      ( cfg_aer_ecrc_check_en ),
    .cfg_aer_ecrc_gen_en                        ( cfg_aer_ecrc_gen_en ),
    .cfg_aer_rooterr_corr_err_reporting_en      ( cfg_aer_rooterr_corr_err_reporting_en ),
    .cfg_aer_rooterr_non_fatal_err_reporting_en ( cfg_aer_rooterr_non_fatal_err_reporting_en ),
    .cfg_aer_rooterr_fatal_err_reporting_en     ( cfg_aer_rooterr_fatal_err_reporting_en ),
    .cfg_aer_rooterr_corr_err_received          ( cfg_aer_rooterr_corr_err_received ),
    .cfg_aer_rooterr_non_fatal_err_received     ( cfg_aer_rooterr_non_fatal_err_received ),
    .cfg_aer_rooterr_fatal_err_received         ( cfg_aer_rooterr_fatal_err_received ),
    .cfg_aer_interrupt_msgnum                   ( cfg_aer_interrupt_msgnum ),
    .cfg_transaction                            ( ),
    .cfg_transaction_addr                       ( ),
    .cfg_transaction_type                       ( ),
    .cfg_vc_tcvc_map                            ( cfg_vc_tcvc_map ),
    .cfg_mgmt_byte_en_n                         ( ~cfg_mgmt_byte_en ),
    .cfg_mgmt_di                                ( cfg_mgmt_di ),
    .cfg_dsn                                    ( cfg_dsn ),
    .cfg_mgmt_dwaddr                            ( cfg_mgmt_dwaddr ),
    .cfg_err_acs_n                              ( 1'b1 ),
    .cfg_err_cor_n                              ( ~cfg_err_cor ),
    .cfg_err_cpl_abort_n                        ( ~cfg_err_cpl_abort ),
    .cfg_err_cpl_timeout_n                      ( ~cfg_err_cpl_timeout ),
    .cfg_err_cpl_unexpect_n                     ( ~cfg_err_cpl_unexpect ),
    .cfg_err_ecrc_n                             ( ~cfg_err_ecrc ),
    .cfg_err_locked_n                           ( ~cfg_err_locked ),
    .cfg_err_posted_n                           ( ~cfg_err_posted ),
    .cfg_err_tlp_cpl_header                     ( cfg_err_tlp_cpl_header ),
    .cfg_err_ur_n                               ( ~cfg_err_ur ),
    .cfg_err_malformed_n                        ( ~cfg_err_malformed ),
    .cfg_err_poisoned_n                         ( ~cfg_err_poisoned ),
    .cfg_err_atomic_egress_blocked_n            ( ~cfg_err_atomic_egress_blocked ),
    .cfg_err_mc_blocked_n                       ( ~cfg_err_mc_blocked ),
    .cfg_err_internal_uncor_n                   ( ~cfg_err_internal_uncor ),
    .cfg_err_internal_cor_n                     ( ~cfg_err_internal_cor ),
    .cfg_err_norecovery_n                       ( ~cfg_err_norecovery ),

    .cfg_interrupt_assert_n                     ( ~cfg_interrupt_assert ),
    .cfg_interrupt_di                           ( cfg_interrupt_di ),
    .cfg_interrupt_n                            ( ~cfg_interrupt ),
    .cfg_interrupt_stat_n                       ( ~cfg_interrupt_stat ),
    .cfg_bus_number                             ( cfg_bus_number ),
    .cfg_device_number                          ( cfg_device_number ),
    .cfg_function_number                        ( cfg_function_number ),
    .cfg_ds_bus_number                          ( cfg_ds_bus_number ),
    .cfg_ds_device_number                       ( cfg_ds_device_number ),
    .cfg_ds_function_number                     ( cfg_ds_function_number ),
    .cfg_pm_send_pme_to_n                       ( 1'b1 ),
    .cfg_pm_wake_n                              ( ~cfg_pm_wake ),
    .cfg_pm_halt_aspm_l0s_n                     ( ~cfg_pm_halt_aspm_l0s ),
    .cfg_pm_halt_aspm_l1_n                      ( ~cfg_pm_halt_aspm_l1 ),
    .cfg_pm_force_state_en_n                    ( ~cfg_pm_force_state_en),
    .cfg_pm_force_state                         ( cfg_pm_force_state ),
    .cfg_force_mps                              ( 3'b0 ),
    .cfg_force_common_clock_off                 ( 1'b0 ),
    .cfg_force_extended_sync_on                 ( 1'b0 ),
    .cfg_port_number                            ( 8'b0 ),
    .cfg_mgmt_rd_en_n                           ( ~cfg_mgmt_rd_en ),
    .cfg_trn_pending                            ( cfg_trn_pending ),
    .cfg_mgmt_wr_en_n                           ( ~cfg_mgmt_wr_en ),
    .cfg_mgmt_wr_readonly_n                     ( ~cfg_mgmt_wr_readonly ),
    .cfg_mgmt_wr_rw1c_as_rw_n                   ( ~cfg_mgmt_wr_rw1c_as_rw ),

    .pl_initial_link_width                      ( pl_initial_link_width ),
    .pl_lane_reversal_mode                      ( pl_lane_reversal_mode ),
    .pl_link_gen2_cap                           ( pl_link_gen2_cap ),
    .pl_link_partner_gen2_supported             ( pl_link_partner_gen2_supported ),
    .pl_link_upcfg_cap                          ( pl_link_upcfg_cap ),
    .pl_phy_lnk_up                              ( pl_phy_lnk_up_wire ),
    .pl_received_hot_rst                        ( pl_received_hot_rst_wire ),
    .pl_rx_pm_state                             ( pl_rx_pm_state ),
    .pl_sel_lnk_rate                            ( pl_sel_lnk_rate ),
    .pl_sel_lnk_width                           ( pl_sel_lnk_width ),
    .pl_tx_pm_state                             ( pl_tx_pm_state ),
    .pl_directed_link_auton                     ( pl_directed_link_auton ),
    .pl_directed_link_change                    ( pl_directed_link_change ),
    .pl_directed_link_speed                     ( pl_directed_link_speed ),
    .pl_directed_link_width                     ( pl_directed_link_width ),
    .pl_downstream_deemph_source                ( pl_downstream_deemph_source ),
    .pl_upstream_prefer_deemph                  ( pl_upstream_prefer_deemph ),
    .pl_transmit_hot_rst                        ( pl_transmit_hot_rst ),
    .pl_directed_ltssm_new_vld                  ( 1'b0 ),
    .pl_directed_ltssm_new                      ( 6'b0 ),
    .pl_directed_ltssm_stall                    ( 1'b0 ),
    .pl_directed_change_done                    ( pl_directed_change_done ),

    .dbg_sclr_a                                 ( ),
    .dbg_sclr_b                                 ( ),
    .dbg_sclr_c                                 ( ),
    .dbg_sclr_d                                 ( ),
    .dbg_sclr_e                                 ( ),
    .dbg_sclr_f                                 ( ),
    .dbg_sclr_g                                 ( ),
    .dbg_sclr_h                                 ( ),
    .dbg_sclr_i                                 ( ),
    .dbg_sclr_j                                 ( ),
    .dbg_sclr_k                                 ( ),

    .dbg_vec_a                                  ( ),
    .dbg_vec_b                                  ( ),
    .dbg_vec_c                                  ( ),
    .pl_dbg_vec                                 ( ),
    .trn_rdllp_data                             ( ),
    .trn_rdllp_src_rdy                          ( ),
    .dbg_mode                                   ( ),
    .dbg_sub_mode                               ( ),
    .pl_dbg_mode                                ( ),

    .drp_clk                                    ( 1'b0 ),
    .drp_do                                     (  ),
    .drp_rdy                                    (  ),
    .drp_addr                                   ( 9'b0 ),
    .drp_en                                     ( 1'b0 ),
    .drp_di                                     ( 16'b0 ),
    .drp_we                                     ( 1'b0 ),

    // Pipe Interface

.pipe_clk                                   ( pipe_clk      ),
.user_clk                                   ( user_clk      ),
.user_clk2                                  ( user_clk2      ),
.phy_rdy_n                                  ( ~phy_rdy      ),

.pl_ltssm_state                             ( pl_ltssm_state_int ),
.pipe_tx_rcvr_det_gt                        ( pipe_tx_rcvr_det_gt    ),
.pipe_tx_rate_gt                            ( common_commands_out[1]     ),
.pipe_tx_deemph_gt                          ( common_commands_out[3]     ),
.pipe_tx_margin_gt                          ( common_commands_out[6:4]  ),


.pipe_tx0_data_gt                           ( pipe_tx_0_sigs[15: 0]      ), 
.pipe_tx0_char_is_k_gt                      ( pipe_tx_0_sigs[17:16]      ),
.pipe_rx0_polarity_gt                       ( pipe_tx_0_sigs[20]         ),
.pipe_tx0_compliance_gt                     ( pipe_tx_0_sigs[19]         ),
.pipe_tx0_elec_idle_gt                      ( pipe_tx_0_sigs[18]         ),
.pipe_tx0_powerdown_gt                      ( pipe_tx_0_sigs[22:21]      ),

.pipe_tx1_data_gt                           ( pipe_tx_1_sigs[15: 0]      ), 
.pipe_tx1_char_is_k_gt                      ( pipe_tx_1_sigs[17:16]      ),
.pipe_rx1_polarity_gt                       ( pipe_tx_1_sigs[20]         ),
.pipe_tx1_compliance_gt                     ( pipe_tx_1_sigs[19]         ),
.pipe_tx1_elec_idle_gt                      ( pipe_tx_1_sigs[18]         ),
.pipe_tx1_powerdown_gt                      ( pipe_tx_1_sigs[22:21]      ),

.pipe_tx2_data_gt                           ( pipe_tx_2_sigs[15: 0]      ), 
.pipe_tx2_char_is_k_gt                      ( pipe_tx_2_sigs[17:16]      ),
.pipe_rx2_polarity_gt                       ( pipe_tx_2_sigs[20]         ),
.pipe_tx2_compliance_gt                     ( pipe_tx_2_sigs[19]         ),
.pipe_tx2_elec_idle_gt                      ( pipe_tx_2_sigs[18]         ),
.pipe_tx2_powerdown_gt                      ( pipe_tx_2_sigs[22:21]      ),

.pipe_tx3_data_gt                           ( pipe_tx_3_sigs[15: 0]      ), 
.pipe_tx3_char_is_k_gt                      ( pipe_tx_3_sigs[17:16]      ),
.pipe_rx3_polarity_gt                       ( pipe_tx_3_sigs[20]         ),
.pipe_tx3_compliance_gt                     ( pipe_tx_3_sigs[19]         ),
.pipe_tx3_elec_idle_gt                      ( pipe_tx_3_sigs[18]         ),
.pipe_tx3_powerdown_gt                      ( pipe_tx_3_sigs[22:21]      ),

.pipe_tx4_data_gt                           ( pipe_tx_4_sigs[15: 0]      ),
.pipe_tx4_char_is_k_gt                      ( pipe_tx_4_sigs[17:16]      ),
.pipe_rx4_polarity_gt                       ( pipe_tx_4_sigs[20]         ),
.pipe_tx4_compliance_gt                     ( pipe_tx_4_sigs[19]         ),
.pipe_tx4_elec_idle_gt                      ( pipe_tx_4_sigs[18]         ),
.pipe_tx4_powerdown_gt                      ( pipe_tx_4_sigs[22:21]      ),

.pipe_tx5_data_gt                           ( pipe_tx_5_sigs[15: 0]      ),
.pipe_tx5_char_is_k_gt                      ( pipe_tx_5_sigs[17:16]      ),
.pipe_rx5_polarity_gt                       ( pipe_tx_5_sigs[20]         ),
.pipe_tx5_compliance_gt                     ( pipe_tx_5_sigs[19]         ),
.pipe_tx5_elec_idle_gt                      ( pipe_tx_5_sigs[18]         ),
.pipe_tx5_powerdown_gt                      ( pipe_tx_5_sigs[22:21]      ),

.pipe_tx6_data_gt                           ( pipe_tx_6_sigs[15: 0]      ),
.pipe_tx6_char_is_k_gt                      ( pipe_tx_6_sigs[17:16]      ),
.pipe_rx6_polarity_gt                       ( pipe_tx_6_sigs[20]         ),
.pipe_tx6_compliance_gt                     ( pipe_tx_6_sigs[19]         ),
.pipe_tx6_elec_idle_gt                      ( pipe_tx_6_sigs[18]         ),
.pipe_tx6_powerdown_gt                      ( pipe_tx_6_sigs[22:21]      ),

.pipe_tx7_data_gt                           ( pipe_tx_7_sigs[15: 0]      ),
.pipe_tx7_char_is_k_gt                      ( pipe_tx_7_sigs[17:16]      ),
.pipe_rx7_polarity_gt                       ( pipe_tx_7_sigs[20]         ),
.pipe_tx7_compliance_gt                     ( pipe_tx_7_sigs[19]         ),
.pipe_tx7_elec_idle_gt                      ( pipe_tx_7_sigs[18]         ),
.pipe_tx7_powerdown_gt                      ( pipe_tx_7_sigs[22:21]      ),

.pipe_rx0_data_gt                           ( pipe_rx_0_sigs[15: 0]      ),
.pipe_rx0_char_is_k_gt                      ( pipe_rx_0_sigs[17:16]      ),
.pipe_rx0_valid_gt                          (~pipe_rx_0_sigs[18]         ),
.pipe_rx0_chanisaligned_gt                  (~pipe_rx_0_sigs[18]         ),
.pipe_rx0_status_gt                         ( rx_status                  ),
.pipe_rx0_phy_status_gt                     ( phy_status                 ),
.pipe_rx0_elec_idle_gt                      ( pipe_rx_0_sigs[18]         ),

.pipe_rx1_data_gt                           ( pipe_rx_1_sigs[15: 0]      ),
.pipe_rx1_char_is_k_gt                      ( pipe_rx_1_sigs[17:16]      ),
.pipe_rx1_valid_gt                          (~pipe_rx_1_sigs[18]         ),
.pipe_rx1_chanisaligned_gt                  (~pipe_rx_1_sigs[18]         ),
.pipe_rx1_status_gt                         ( rx_status              ),
.pipe_rx1_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH >= 2 )? phy_status : 1'b0   ),
.pipe_rx1_elec_idle_gt                      ( pipe_rx_1_sigs[18]         ),

.pipe_rx2_data_gt                           ( pipe_rx_2_sigs[15: 0]      ),
.pipe_rx2_char_is_k_gt                      ( pipe_rx_2_sigs[17:16]      ),
.pipe_rx2_valid_gt                          (~pipe_rx_2_sigs[18]         ),
.pipe_rx2_chanisaligned_gt                  (~pipe_rx_2_sigs[18]         ),
.pipe_rx2_status_gt                         ( rx_status                  ),
.pipe_rx2_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0          ),
.pipe_rx2_elec_idle_gt                      ( pipe_rx_2_sigs[18]         ),

.pipe_rx3_data_gt                           ( pipe_rx_3_sigs[15: 0]      ),
.pipe_rx3_char_is_k_gt                      ( pipe_rx_3_sigs[17:16]      ),
.pipe_rx3_valid_gt                          (~pipe_rx_3_sigs[18]         ),
.pipe_rx3_chanisaligned_gt                  (~pipe_rx_3_sigs[18]         ),
.pipe_rx3_status_gt                         ( rx_status                  ),
.pipe_rx3_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0          ),
.pipe_rx3_elec_idle_gt                      ( pipe_rx_3_sigs[18]         ),

.pipe_rx4_data_gt                           ( pipe_rx_4_sigs[15: 0]      ),
.pipe_rx4_char_is_k_gt                      ( pipe_rx_4_sigs[17:16]      ),
.pipe_rx4_valid_gt                          (~pipe_rx_4_sigs[18]         ),
.pipe_rx4_chanisaligned_gt                  (~pipe_rx_4_sigs[18]         ),
.pipe_rx4_status_gt                         ( rx_status     ),
.pipe_rx4_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH == 8 )? phy_status : 1'b0        ),
.pipe_rx4_elec_idle_gt                      ( pipe_rx_4_sigs[18]         ),

.pipe_rx5_data_gt                           ( pipe_rx_5_sigs[15: 0]      ),
.pipe_rx5_char_is_k_gt                      ( pipe_rx_5_sigs[17:16]      ),
.pipe_rx5_valid_gt                          (~pipe_rx_5_sigs[18]         ),
.pipe_rx5_chanisaligned_gt                  (~pipe_rx_5_sigs[18]         ),
.pipe_rx5_status_gt                         ( rx_status      ),
.pipe_rx5_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH == 8 )? phy_status : 1'b0        ),
.pipe_rx5_elec_idle_gt                      ( pipe_rx_5_sigs[18]         ),

.pipe_rx6_data_gt                           ( pipe_rx_6_sigs[15: 0]      ),
.pipe_rx6_char_is_k_gt                      ( pipe_rx_6_sigs[17:16]      ),
.pipe_rx6_valid_gt                          (~pipe_rx_6_sigs[18]         ),
.pipe_rx6_chanisaligned_gt                  (~pipe_rx_6_sigs[18]         ),
.pipe_rx6_status_gt                         ( rx_status      ),
.pipe_rx6_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH == 8 )? phy_status : 1'b0      ),
.pipe_rx6_elec_idle_gt                      ( pipe_rx_6_sigs[18]         ),

.pipe_rx7_data_gt                           ( pipe_rx_7_sigs[15: 0]      ),
.pipe_rx7_char_is_k_gt                      ( pipe_rx_7_sigs[17:16]      ),
.pipe_rx7_valid_gt                          (~pipe_rx_7_sigs[18]         ),
.pipe_rx7_chanisaligned_gt                  (~pipe_rx_7_sigs[18]         ),
.pipe_rx7_status_gt                         ( rx_status     ),
.pipe_rx7_phy_status_gt                     ( (LINK_CAP_MAX_LINK_WIDTH == 8 )? phy_status : 1'b0         ),
.pipe_rx7_elec_idle_gt                      ( pipe_rx_7_sigs[18]         )

);
// Pipe mode tie-offs
assign common_commands_out[0] = pipe_clk;
assign common_commands_out[2] = pipe_tx_rcvr_det_gt;
assign common_commands_out[11:7] = 5'b0;  

end
endgenerate

generate if (EXT_PIPE_SIM == "FALSE")
begin

  //------------------------------------------------------------------------------------------------------------------//
  // **** V7/K7/A7 GTX Wrapper ****                                                                                   //
  //   The 7-Series GTX Wrapper includes the following:                                                               //
  //     1) Virtex-7 GTX                                                                                              //
  //     2) Kintex-7 GTX                                                                                              //
  //     3) Artix-7  GTP                                                                                              //
  //------------------------------------------------------------------------------------------------------------------//
model_ap2_tst_gt_top #(
    .LINK_CAP_MAX_LINK_WIDTH       ( LINK_CAP_MAX_LINK_WIDTH ),
    .REF_CLK_FREQ                  ( REF_CLK_FREQ ),
    .USER_CLK_FREQ                 ( USER_CLK_FREQ ),
    .USER_CLK2_DIV2                ( USER_CLK2_DIV2 ),
    .PL_FAST_TRAIN                 ( PL_FAST_TRAIN ),
    .PCIE_EXT_CLK                  ( PCIE_EXT_CLK ),
    .PCIE_USE_MODE                 ( PCIE_USE_MODE ),
    .PCIE_GT_DEVICE                ( PCIE_GT_DEVICE ),
    .PCIE_PLL_SEL                  ( PCIE_PLL_SEL ),
    .PCIE_ASYNC_EN                 ( PCIE_ASYNC_EN ),
    .PCIE_TXBUF_EN                 ( PCIE_TXBUF_EN ),
    .PCIE_CHAN_BOND                ( PCIE_CHAN_BOND )
  ) model_ap2_tst_gt_top_i (
    // pl ltssm
    .pl_ltssm_state                ( pl_ltssm_state_int ),

    // Pipe Common Signals
    .pipe_tx_rcvr_det              ( pipe_tx_rcvr_det_gt  ),
    .pipe_tx_reset                 ( 1'b0                 ),
    .pipe_tx_rate                  ( pipe_tx_rate_gt      ),
    .pipe_tx_deemph                ( pipe_tx_deemph_gt    ),
    .pipe_tx_margin                ( pipe_tx_margin_gt    ),
    .pipe_tx_swing                 ( 1'b0                 ),

    // Pipe Per-Lane Signals - Lane 0
    .pipe_rx0_char_is_k            ( pipe_rx0_char_is_k_gt),
    .pipe_rx0_data                 ( pipe_rx0_data_gt     ),
    .pipe_rx0_valid                ( pipe_rx0_valid_gt    ),
    .pipe_rx0_chanisaligned        ( pipe_rx0_chanisaligned_gt   ),
    .pipe_rx0_status               ( pipe_rx0_status_gt      ),
    .pipe_rx0_phy_status           ( pipe_rx0_phy_status_gt  ),
    .pipe_rx0_elec_idle            ( pipe_rx0_elec_idle_gt   ),
    .pipe_rx0_polarity             ( pipe_rx0_polarity_gt    ),
    .pipe_tx0_compliance           ( pipe_tx0_compliance_gt  ),
    .pipe_tx0_char_is_k            ( pipe_tx0_char_is_k_gt   ),
    .pipe_tx0_data                 ( pipe_tx0_data_gt        ),
    .pipe_tx0_elec_idle            ( pipe_tx0_elec_idle_gt   ),
    .pipe_tx0_powerdown            ( pipe_tx0_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 1

    .pipe_rx1_char_is_k            ( pipe_rx1_char_is_k_gt),
    .pipe_rx1_data                 ( pipe_rx1_data_gt     ),
    .pipe_rx1_valid                ( pipe_rx1_valid_gt    ),
    .pipe_rx1_chanisaligned        ( pipe_rx1_chanisaligned_gt   ),
    .pipe_rx1_status               ( pipe_rx1_status_gt      ),
    .pipe_rx1_phy_status           ( pipe_rx1_phy_status_gt  ),
    .pipe_rx1_elec_idle            ( pipe_rx1_elec_idle_gt   ),
    .pipe_rx1_polarity             ( pipe_rx1_polarity_gt    ),
    .pipe_tx1_compliance           ( pipe_tx1_compliance_gt  ),
    .pipe_tx1_char_is_k            ( pipe_tx1_char_is_k_gt   ),
    .pipe_tx1_data                 ( pipe_tx1_data_gt        ),
    .pipe_tx1_elec_idle            ( pipe_tx1_elec_idle_gt   ),
    .pipe_tx1_powerdown            ( pipe_tx1_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 2

    .pipe_rx2_char_is_k            ( pipe_rx2_char_is_k_gt),
    .pipe_rx2_data                 ( pipe_rx2_data_gt     ),
    .pipe_rx2_valid                ( pipe_rx2_valid_gt    ),
    .pipe_rx2_chanisaligned        ( pipe_rx2_chanisaligned_gt   ),
    .pipe_rx2_status               ( pipe_rx2_status_gt      ),
    .pipe_rx2_phy_status           ( pipe_rx2_phy_status_gt  ),
    .pipe_rx2_elec_idle            ( pipe_rx2_elec_idle_gt   ),
    .pipe_rx2_polarity             ( pipe_rx2_polarity_gt    ),
    .pipe_tx2_compliance           ( pipe_tx2_compliance_gt  ),
    .pipe_tx2_char_is_k            ( pipe_tx2_char_is_k_gt   ),
    .pipe_tx2_data                 ( pipe_tx2_data_gt        ),
    .pipe_tx2_elec_idle            ( pipe_tx2_elec_idle_gt   ),
    .pipe_tx2_powerdown            ( pipe_tx2_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 3

    .pipe_rx3_char_is_k            ( pipe_rx3_char_is_k_gt),
    .pipe_rx3_data                 ( pipe_rx3_data_gt     ),
    .pipe_rx3_valid                ( pipe_rx3_valid_gt    ),
    .pipe_rx3_chanisaligned        ( pipe_rx3_chanisaligned_gt   ),
    .pipe_rx3_status               ( pipe_rx3_status_gt      ),
    .pipe_rx3_phy_status           ( pipe_rx3_phy_status_gt  ),
    .pipe_rx3_elec_idle            ( pipe_rx3_elec_idle_gt   ),
    .pipe_rx3_polarity             ( pipe_rx3_polarity_gt    ),
    .pipe_tx3_compliance           ( pipe_tx3_compliance_gt  ),
    .pipe_tx3_char_is_k            ( pipe_tx3_char_is_k_gt   ),
    .pipe_tx3_data                 ( pipe_tx3_data_gt        ),
    .pipe_tx3_elec_idle            ( pipe_tx3_elec_idle_gt   ),
    .pipe_tx3_powerdown            ( pipe_tx3_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 4

    .pipe_rx4_char_is_k            ( pipe_rx4_char_is_k_gt),
    .pipe_rx4_data                 ( pipe_rx4_data_gt     ),
    .pipe_rx4_valid                ( pipe_rx4_valid_gt    ),
    .pipe_rx4_chanisaligned        ( pipe_rx4_chanisaligned_gt   ),
    .pipe_rx4_status               ( pipe_rx4_status_gt      ),
    .pipe_rx4_phy_status           ( pipe_rx4_phy_status_gt  ),
    .pipe_rx4_elec_idle            ( pipe_rx4_elec_idle_gt   ),
    .pipe_rx4_polarity             ( pipe_rx4_polarity_gt    ),
    .pipe_tx4_compliance           ( pipe_tx4_compliance_gt  ),
    .pipe_tx4_char_is_k            ( pipe_tx4_char_is_k_gt   ),
    .pipe_tx4_data                 ( pipe_tx4_data_gt        ),
    .pipe_tx4_elec_idle            ( pipe_tx4_elec_idle_gt   ),
    .pipe_tx4_powerdown            ( pipe_tx4_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 5

    .pipe_rx5_char_is_k            ( pipe_rx5_char_is_k_gt),
    .pipe_rx5_data                 ( pipe_rx5_data_gt     ),
    .pipe_rx5_valid                ( pipe_rx5_valid_gt    ),
    .pipe_rx5_chanisaligned        ( pipe_rx5_chanisaligned_gt   ),
    .pipe_rx5_status               ( pipe_rx5_status_gt      ),
    .pipe_rx5_phy_status           ( pipe_rx5_phy_status_gt  ),
    .pipe_rx5_elec_idle            ( pipe_rx5_elec_idle_gt   ),
    .pipe_rx5_polarity             ( pipe_rx5_polarity_gt    ),
    .pipe_tx5_compliance           ( pipe_tx5_compliance_gt  ),
    .pipe_tx5_char_is_k            ( pipe_tx5_char_is_k_gt   ),
    .pipe_tx5_data                 ( pipe_tx5_data_gt        ),
    .pipe_tx5_elec_idle            ( pipe_tx5_elec_idle_gt   ),
    .pipe_tx5_powerdown            ( pipe_tx5_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 6

    .pipe_rx6_char_is_k            ( pipe_rx6_char_is_k_gt),
    .pipe_rx6_data                 ( pipe_rx6_data_gt     ),
    .pipe_rx6_valid                ( pipe_rx6_valid_gt    ),
    .pipe_rx6_chanisaligned        ( pipe_rx6_chanisaligned_gt   ),
    .pipe_rx6_status               ( pipe_rx6_status_gt      ),
    .pipe_rx6_phy_status           ( pipe_rx6_phy_status_gt  ),
    .pipe_rx6_elec_idle            ( pipe_rx6_elec_idle_gt   ),
    .pipe_rx6_polarity             ( pipe_rx6_polarity_gt    ),
    .pipe_tx6_compliance           ( pipe_tx6_compliance_gt  ),
    .pipe_tx6_char_is_k            ( pipe_tx6_char_is_k_gt   ),
    .pipe_tx6_data                 ( pipe_tx6_data_gt        ),
    .pipe_tx6_elec_idle            ( pipe_tx6_elec_idle_gt   ),
    .pipe_tx6_powerdown            ( pipe_tx6_powerdown_gt   ),

    // Pipe Per-Lane Signals - Lane 7

    .pipe_rx7_char_is_k            ( pipe_rx7_char_is_k_gt),
    .pipe_rx7_data                 ( pipe_rx7_data_gt     ),
    .pipe_rx7_valid                ( pipe_rx7_valid_gt    ),
    .pipe_rx7_chanisaligned        ( pipe_rx7_chanisaligned_gt   ),
    .pipe_rx7_status               ( pipe_rx7_status_gt      ),
    .pipe_rx7_phy_status           ( pipe_rx7_phy_status_gt  ),
    .pipe_rx7_elec_idle            ( pipe_rx7_elec_idle_gt   ),
    .pipe_rx7_polarity             ( pipe_rx7_polarity_gt    ),
    .pipe_tx7_compliance           ( pipe_tx7_compliance_gt  ),
    .pipe_tx7_char_is_k            ( pipe_tx7_char_is_k_gt   ),
    .pipe_tx7_data                 ( pipe_tx7_data_gt        ),
    .pipe_tx7_elec_idle            ( pipe_tx7_elec_idle_gt   ),
    .pipe_tx7_powerdown            ( pipe_tx7_powerdown_gt   ),

    // PCI Express Signals
    .pci_exp_txn                   ( pci_exp_txn          ),
    .pci_exp_txp                   ( pci_exp_txp          ),
    .pci_exp_rxn                   ( pci_exp_rxn          ),
    .pci_exp_rxp                   ( pci_exp_rxp          ),

    // Non PIPE Signals
    .sys_clk                       ( sys_clk             ),
    .sys_rst_n                     ( sys_rst_n           ),
    .PIPE_MMCM_RST_N               ( pipe_mmcm_rst_n     ),        // Async      | Async
    .pipe_clk                      ( pipe_clk            ),

    .user_clk                      ( user_clk            ),
    .user_clk2                     ( user_clk2           ),
    .phy_rdy_n                     ( phy_rdy_n           ),

    .PIPE_PCLK_IN                  ( pipe_pclk_in ),
    .PIPE_RXUSRCLK_IN              ( pipe_rxusrclk_in ),
    .PIPE_RXOUTCLK_IN              ( pipe_rxoutclk_in ),
    .PIPE_DCLK_IN                  ( pipe_dclk_in ),
    .PIPE_USERCLK1_IN              ( pipe_userclk1_in ),
    .PIPE_USERCLK2_IN              ( pipe_userclk2_in ),
    .PIPE_OOBCLK_IN                ( pipe_oobclk_in ),
    .PIPE_MMCM_LOCK_IN             ( pipe_mmcm_lock_in ),

    .PIPE_TXOUTCLK_OUT             ( pipe_txoutclk_out ),
    .PIPE_RXOUTCLK_OUT             ( pipe_rxoutclk_out ),
    .PIPE_PCLK_SEL_OUT             ( pipe_pclk_sel_out ),
    .PIPE_GEN3_OUT                 ( pipe_gen3_out ),

     //-----------External GT COMMON Ports-----------------------------------

    .qpll_drp_crscode               (  ),
    .qpll_drp_fsm                   (  ),
    .qpll_drp_done                  (  ), 
    .qpll_drp_reset                 (  ),
    .qpll_qplllock                  (  ),
    .qpll_qplloutclk                (  ),
    .qpll_qplloutrefclk             (  ) ,
    .qpll_qplld                     ( qpll_qplld ),
    .qpll_qpllreset                 (  ),
    .qpll_drp_clk                   ( qpll_drp_clk ),
    .qpll_drp_rst_n                 ( qpll_drp_rst_n ),
    .qpll_drp_ovrd                  ( qpll_drp_ovrd ),
    .qpll_drp_gen3                  ( qpll_drp_gen3),
    .qpll_drp_start                 ( qpll_drp_start ),
 
    //TRANSCEIVER DEBUG EOU
    .ext_ch_gt_drpclk               (  ),
    .ext_ch_gt_drpaddr              (36'd0 ),
    .ext_ch_gt_drpen                (4'd0),
    .ext_ch_gt_drpdi                (64'd0),
    .ext_ch_gt_drpwe                (4'd0  ),
    .ext_ch_gt_drpdo                (  ),
    .ext_ch_gt_drprdy               (  ),

    //---------- PRBS/Loopback Ports -----------------------
    .PIPE_TXPRBSSEL                (  ), 
    .PIPE_RXPRBSSEL                (  ), 
    .PIPE_TXPRBSFORCEERR           (  ), 
    .PIPE_RXPRBSCNTRESET           (  ), 
    .PIPE_LOOPBACK                 (  ), 

    .PIPE_RXPRBSERR                ( ),

     //---------- Transceiver Debug FSM Ports ---------------------------------
    .PIPE_RST_FSM                  ( ),
    .PIPE_QRST_FSM                 ( ),
    .PIPE_RATE_FSM                 ( ),
    .PIPE_SYNC_FSM_TX              ( ),
    .PIPE_SYNC_FSM_RX              ( ),
    .PIPE_DRP_FSM                  ( ),

    .PIPE_RST_IDLE                 ( pipe_rst_idle ),
    .PIPE_QRST_IDLE                ( pipe_qrst_idle ),
    .PIPE_RATE_IDLE                ( pipe_rate_idle ),
    .PIPE_EYESCANDATAERROR         ( ),
    .PIPE_RXSTATUS                 ( ), 
    .PIPE_DMONITOROUT              ( ),

    .PIPE_CPLL_LOCK                ( ), 
    .PIPE_QPLL_LOCK                ( ), 
    .PIPE_RXPMARESETDONE           ( ),       
    .PIPE_RXBUFSTATUS              ( ),      
    .PIPE_TXPHALIGNDONE            ( ),      
    .PIPE_TXPHINITDONE             ( ),      
    .PIPE_TXDLYSRESETDONE          ( ),     
    .PIPE_RXPHALIGNDONE            ( ),     
    .PIPE_RXDLYSRESETDONE          ( ),      
    .PIPE_RXSYNCDONE               ( ),   
    .PIPE_RXDISPERR                ( ),  
    .PIPE_RXNOTINTABLE             ( ),    
    .PIPE_RXCOMMADET               ( ),    
    //---------- JTAG Ports --------------------------------
    .PIPE_JTAG_RDY                 ( ),

   //---------- Debug Ports -------------------------------
    .PIPE_DEBUG_0                  ( ),
    .PIPE_DEBUG_1                  ( ),
    .PIPE_DEBUG_2                  ( ),
    .PIPE_DEBUG_3                  ( ),
    .PIPE_DEBUG_4                  ( ),
    .PIPE_DEBUG_5                  ( ),
    .PIPE_DEBUG_6                  ( ),
    .PIPE_DEBUG_7                  ( ),
    .PIPE_DEBUG_8                  ( ),
    .PIPE_DEBUG_9                  ( ),
    .PIPE_DEBUG                    ( ),
    .INT_PCLK_SEL_SLAVE(),
    .INT_QPLLOUTREFCLK_OUT(),
    .INT_QPLLOUTCLK_OUT(),
    .INT_QPLLLOCK_OUT(),
    .INT_MMCM_LOCK_OUT(),
    .INT_OOBCLK_OUT(),
    .INT_USERCLK2_OUT(),
    .INT_USERCLK1_OUT(),
    .INT_DCLK_OUT(),
    .INT_RXOUTCLK_OUT(),
    .INT_RXUSRCLK_OUT(),
    .INT_PCLK_OUT_SLAVE()
  );
end
endgenerate

//  assign  common_commands_out = 12'b0;  
//  assign  pipe_tx_0_sigs      = 25'b0;   
//  assign  pipe_tx_1_sigs      = 25'b0; 
//  assign  pipe_tx_2_sigs      = 25'b0; 
//  assign  pipe_tx_3_sigs      = 25'b0; 
//  assign  pipe_tx_4_sigs      = 25'b0; 
//  assign  pipe_tx_5_sigs      = 25'b0; 
//  assign  pipe_tx_6_sigs      = 25'b0; 
//  assign  pipe_tx_7_sigs      = 25'b0; 

endmodule


`timescale 1ns/1ps
module model_ap2_tst_pcie_top # (
  // PCIE_2_1 params
  parameter        PIPE_PIPELINE_STAGES = 0,                // 0 - 0 stages, 1 - 1 stage, 2 - 2 stages
  parameter [11:0] AER_BASE_PTR = 12'h140,
  parameter        AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter        DEV_CAP_ROLE_BASED_ERROR = "TRUE",
  parameter        LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE",
  parameter        AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [15:0] AER_CAP_ID = 16'h0001,
  parameter        AER_CAP_MULTIHEADER = "FALSE",
  parameter [11:0] AER_CAP_NEXTPTR = 12'h178,
  parameter        AER_CAP_ON = "FALSE",
  parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000,
  parameter        AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE",
  parameter [3:0]  AER_CAP_VERSION = 4'h1,
  parameter        ALLOW_X8_GEN2 = "FALSE",
  parameter [31:0] BAR0 = 32'hFFFFFF00,
  parameter [31:0] BAR1 = 32'hFFFF0000,
  parameter [31:0] BAR2 = 32'hFFFF000C,
  parameter [31:0] BAR3 = 32'hFFFFFFFF,
  parameter [31:0] BAR4 = 32'h00000000,
  parameter [31:0] BAR5 = 32'h00000000,
  parameter        C_DATA_WIDTH = 64,
  parameter        REM_WIDTH = (C_DATA_WIDTH == 128) ? 2 : 1,
  parameter        KEEP_WIDTH = C_DATA_WIDTH / 8,
  parameter [7:0]  CAPABILITIES_PTR = 8'h40,
  parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000,
  parameter [23:0] CLASS_CODE = 24'h000000,
  parameter        CFG_ECRC_ERR_CPLSTAT = 0,
  parameter        CMD_INTX_IMPLEMENTED = "TRUE",
  parameter        CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE",
  parameter [3:0]  CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0,
  parameter [6:0]  CRM_MODULE_RSTS = 7'h00,
  parameter        DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE",
  parameter [1:0]  DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0,
  parameter        DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE",
  parameter [1:0]  DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0,
  parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE",
  parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE",
  parameter        integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0,
  parameter        integer DEV_CAP_ENDPOINT_L1_LATENCY = 0,
  parameter        DEV_CAP_EXT_TAG_SUPPORTED = "TRUE",
  parameter        DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE",
  parameter        integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2,
  parameter        integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0,
  parameter        integer DEV_CAP_RSVD_14_12 = 0,
  parameter        integer DEV_CAP_RSVD_17_16 = 0,
  parameter        integer DEV_CAP_RSVD_31_29 = 0,
  parameter        DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE",
  parameter        DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE",
  parameter        DISABLE_ASPM_L1_TIMER = "FALSE",
  parameter        DISABLE_BAR_FILTERING = "FALSE",
  parameter        DISABLE_ERR_MSG = "FALSE",
  parameter        DISABLE_ID_CHECK = "FALSE",
  parameter        DISABLE_LANE_REVERSAL = "FALSE",
  parameter        DISABLE_LOCKED_FILTER = "FALSE",
  parameter        DISABLE_PPM_FILTER = "FALSE",
  parameter        DISABLE_RX_POISONED_RESP = "FALSE",
  parameter        DISABLE_RX_TC_FILTER = "FALSE",
  parameter        DISABLE_SCRAMBLING = "FALSE",
  parameter [7:0]  DNSTREAM_LINK_NUM = 8'h00,
  parameter [11:0] DSN_BASE_PTR = 12'h100,
  parameter [15:0] DSN_CAP_ID = 16'h0003,
  parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C,
  parameter        DSN_CAP_ON = "TRUE",
  parameter [3:0]  DSN_CAP_VERSION = 4'h1,
  parameter [10:0] ENABLE_MSG_ROUTE = 11'h000,
  parameter        ENABLE_RX_TD_ECRC_TRIM = "FALSE",
  parameter        ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE",
  parameter        ENTER_RVRY_EI_L0 = "TRUE",
  parameter        EXIT_LOOPBACK_ON_EI = "TRUE",
  parameter [31:0] EXPANSION_ROM = 32'hFFFFF001,
  parameter [5:0]  EXT_CFG_CAP_PTR = 6'h3F,
  parameter [9:0]  EXT_CFG_XP_CAP_PTR = 10'h3FF,
  parameter [7:0]  HEADER_TYPE = 8'h00,
  parameter [4:0]  INFER_EI = 5'h00,
  parameter [7:0]  INTERRUPT_PIN = 8'h01,
  parameter        INTERRUPT_STAT_AUTO = "TRUE",
  parameter        IS_SWITCH = "FALSE",
  parameter [9:0]  LAST_CONFIG_DWORD = 10'h3FF,
  parameter        LINK_CAP_ASPM_OPTIONALITY = "TRUE",
  parameter        integer LINK_CAP_ASPM_SUPPORT = 1,
  parameter        LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE",
  parameter        LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE",
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7,
  parameter        LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE",
  parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,
  parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,
  parameter        integer LINK_CAP_RSVD_23 = 0,
  parameter        integer LINK_CONTROL_RCB = 0,
  parameter        LINK_CTRL2_DEEMPHASIS = "FALSE",
  parameter        LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE",
  parameter [3:0]  LINK_CTRL2_TARGET_LINK_SPEED = 4'h2,
  parameter        LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE",
  parameter [14:0] LL_ACK_TIMEOUT = 15'h0000,
  parameter        LL_ACK_TIMEOUT_EN = "FALSE",
  parameter        integer LL_ACK_TIMEOUT_FUNC = 0,
  parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000,
  parameter        LL_REPLAY_TIMEOUT_EN = "FALSE",
  parameter        integer LL_REPLAY_TIMEOUT_FUNC = 0,
  parameter [5:0]  LTSSM_MAX_LINK_WIDTH = 6'h01,
  parameter        MPS_FORCE = "FALSE",
  parameter [7:0]  MSIX_BASE_PTR = 8'h9C,
  parameter [7:0]  MSIX_CAP_ID = 8'h11,
  parameter [7:0]  MSIX_CAP_NEXTPTR = 8'h00,
  parameter        MSIX_CAP_ON = "FALSE",
  parameter        integer MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter        integer MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter [7:0]  MSI_BASE_PTR = 8'h48,
  parameter        MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE",
  parameter [7:0]  MSI_CAP_ID = 8'h05,
  parameter        integer MSI_CAP_MULTIMSGCAP = 0,
  parameter        integer MSI_CAP_MULTIMSG_EXTENSION = 0,
  parameter [7:0]  MSI_CAP_NEXTPTR = 8'h60,
  parameter        MSI_CAP_ON = "FALSE",
  parameter        MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE",
  parameter        integer N_FTS_COMCLK_GEN1 = 255,
  parameter        integer N_FTS_COMCLK_GEN2 = 255,
  parameter        integer N_FTS_GEN1 = 255,
  parameter        integer N_FTS_GEN2 = 255,
  parameter [7:0]  PCIE_BASE_PTR = 8'h60,
  parameter [7:0]  PCIE_CAP_CAPABILITY_ID = 8'h10,
  parameter [3:0]  PCIE_CAP_CAPABILITY_VERSION = 4'h2,
  parameter [3:0]  PCIE_CAP_DEVICE_PORT_TYPE = 4'h0,
  parameter [7:0]  PCIE_CAP_NEXTPTR = 8'h9C,
  parameter        PCIE_CAP_ON = "TRUE",
  parameter        integer PCIE_CAP_RSVD_15_14 = 0,
  parameter        PCIE_CAP_SLOT_IMPLEMENTED = "FALSE",
  parameter        integer PCIE_REVISION = 2,
  parameter        integer PL_AUTO_CONFIG = 0,
  parameter        PL_FAST_TRAIN = "FALSE",
  parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000,
  parameter        PM_ASPML0S_TIMEOUT_EN = "FALSE",
  parameter        integer PM_ASPML0S_TIMEOUT_FUNC = 0,
  parameter        PM_ASPM_FASTEXIT = "FALSE",
  parameter [7:0]  PM_BASE_PTR = 8'h40,
  parameter        integer PM_CAP_AUXCURRENT = 0,
  parameter        PM_CAP_D1SUPPORT = "TRUE",
  parameter        PM_CAP_D2SUPPORT = "TRUE",
  parameter        PM_CAP_DSI = "FALSE",
  parameter [7:0]  PM_CAP_ID = 8'h01,
  parameter [7:0]  PM_CAP_NEXTPTR = 8'h48,
  parameter        PM_CAP_ON = "TRUE",
  parameter [4:0]  PM_CAP_PMESUPPORT = 5'h0F,
  parameter        PM_CAP_PME_CLOCK = "FALSE",
  parameter        integer PM_CAP_RSVD_04 = 0,
  parameter        integer PM_CAP_VERSION = 3,
  parameter        PM_CSR_B2B3 = "FALSE",
  parameter        PM_CSR_BPCCEN = "FALSE",
  parameter        PM_CSR_NOSOFTRST = "TRUE",
  parameter [7:0]  PM_DATA0 = 8'h01,
  parameter [7:0]  PM_DATA1 = 8'h01,
  parameter [7:0]  PM_DATA2 = 8'h01,
  parameter [7:0]  PM_DATA3 = 8'h01,
  parameter [7:0]  PM_DATA4 = 8'h01,
  parameter [7:0]  PM_DATA5 = 8'h01,
  parameter [7:0]  PM_DATA6 = 8'h01,
  parameter [7:0]  PM_DATA7 = 8'h01,
  parameter [1:0]  PM_DATA_SCALE0 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE1 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE2 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE3 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE4 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE5 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE6 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE7 = 2'h1,
  parameter        PM_MF = "FALSE",
  parameter [11:0] RBAR_BASE_PTR = 12'h178,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00,
  parameter [15:0] RBAR_CAP_ID = 16'h0015,
  parameter [2:0]  RBAR_CAP_INDEX0 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX1 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX2 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX3 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX4 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX5 = 3'h0,
  parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000,
  parameter        RBAR_CAP_ON = "FALSE",
  parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000,
  parameter [3:0]  RBAR_CAP_VERSION = 4'h1,
  parameter [2:0]  RBAR_NUM = 3'h1,
  parameter        integer RECRC_CHK = 0,
  parameter        RECRC_CHK_TRIM = "FALSE",
  parameter        ROOT_CAP_CRS_SW_VISIBILITY = "FALSE",
  parameter [1:0]  RP_AUTO_SPD = 2'h1,
  parameter [4:0]  RP_AUTO_SPD_LOOPCNT = 5'h1f,
  parameter        SELECT_DLL_IF = "FALSE",
  parameter        SIM_VERSION = "1.0",
  parameter        SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE",
  parameter        SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE",
  parameter        SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE",
  parameter        SLOT_CAP_HOTPLUG_CAPABLE = "FALSE",
  parameter        SLOT_CAP_HOTPLUG_SURPRISE = "FALSE",
  parameter        SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE",
  parameter        SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE",
  parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000,
  parameter        SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE",
  parameter        SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE",
  parameter        integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0,
  parameter [7:0]  SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00,
  parameter        integer SPARE_BIT0 = 0,
  parameter        integer SPARE_BIT1 = 0,
  parameter        integer SPARE_BIT2 = 0,
  parameter        integer SPARE_BIT3 = 0,
  parameter        integer SPARE_BIT4 = 0,
  parameter        integer SPARE_BIT5 = 0,
  parameter        integer SPARE_BIT6 = 0,
  parameter        integer SPARE_BIT7 = 0,
  parameter        integer SPARE_BIT8 = 0,
  parameter [7:0]  SPARE_BYTE0 = 8'h00,
  parameter [7:0]  SPARE_BYTE1 = 8'h00,
  parameter [7:0]  SPARE_BYTE2 = 8'h00,
  parameter [7:0]  SPARE_BYTE3 = 8'h00,
  parameter [31:0] SPARE_WORD0 = 32'h00000000,
  parameter [31:0] SPARE_WORD1 = 32'h00000000,
  parameter [31:0] SPARE_WORD2 = 32'h00000000,
  parameter [31:0] SPARE_WORD3 = 32'h00000000,
  parameter        SSL_MESSAGE_AUTO = "FALSE",
  parameter        TECRC_EP_INV = "FALSE",
  parameter        TL_RBYPASS = "FALSE",
  parameter        integer TL_RX_RAM_RADDR_LATENCY = 0,
  parameter        integer TL_RX_RAM_RDATA_LATENCY = 2,
  parameter        integer TL_RX_RAM_WRITE_LATENCY = 0,
  parameter        TL_TFC_DISABLE = "FALSE",
  parameter        TL_TX_CHECKS_DISABLE = "FALSE",
  parameter        integer TL_TX_RAM_RADDR_LATENCY = 0,
  parameter        integer TL_TX_RAM_RDATA_LATENCY = 2,
  parameter        integer TL_TX_RAM_WRITE_LATENCY = 0,
  parameter        TRN_DW = "FALSE",
  parameter        TRN_NP_FC = "FALSE",
  parameter        UPCONFIG_CAPABLE = "TRUE",
  parameter        UPSTREAM_FACING = "TRUE",
  parameter        UR_ATOMIC = "TRUE",
  parameter        UR_CFG1 = "TRUE",
  parameter        UR_INV_REQ = "TRUE",
  parameter        UR_PRS_RESPONSE = "TRUE",
  parameter        USER_CLK2_DIV2 = "FALSE",
  parameter        integer USER_CLK_FREQ = 3,
  parameter        USE_RID_PINS = "FALSE",
  parameter        VC0_CPL_INFINITE = "TRUE",
  parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF,
  parameter        integer VC0_TOTAL_CREDITS_CD = 127,
  parameter        integer VC0_TOTAL_CREDITS_CH = 31,
  parameter        integer VC0_TOTAL_CREDITS_NPD = 24,
  parameter        integer VC0_TOTAL_CREDITS_NPH = 12,
  parameter        integer VC0_TOTAL_CREDITS_PD = 288,
  parameter        integer VC0_TOTAL_CREDITS_PH = 32,
  parameter        integer VC0_TX_LASTPACKET = 31,
  parameter [11:0] VC_BASE_PTR = 12'h10C,
  parameter [15:0] VC_CAP_ID = 16'h0002,
  parameter [11:0] VC_CAP_NEXTPTR = 12'h000,
  parameter        VC_CAP_ON = "FALSE",
  parameter        VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE",
  parameter [3:0]  VC_CAP_VERSION = 4'h1,
  parameter [11:0] VSEC_BASE_PTR = 12'h128,
  parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234,
  parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018,
  parameter [3:0]  VSEC_CAP_HDR_REVISION = 4'h1,
  parameter [15:0] VSEC_CAP_ID = 16'h000B,
  parameter        VSEC_CAP_IS_LINK_VISIBLE = "TRUE",
  parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140,
  parameter        VSEC_CAP_ON = "FALSE",
  parameter [3:0]  VSEC_CAP_VERSION = 4'h1
)
(

  // wrapper input
  // Common
  output                                     user_clk_out,
  input                                      user_reset,
  input                                      user_lnk_up,

  output                                     trn_lnk_up,
  output                                     user_rst_n,

  // Tx
  output  [5:0]                              tx_buf_av,
  output                                     tx_err_drop,
  output                                     tx_cfg_req,
  output                                     s_axis_tx_tready,
  input   [C_DATA_WIDTH-1:0]                 s_axis_tx_tdata,
  input   [KEEP_WIDTH-1:0]                   s_axis_tx_tkeep,
  input   [3:0]                              s_axis_tx_tuser,
  input                                      s_axis_tx_tlast,
  input                                      s_axis_tx_tvalid,
  input                                      tx_cfg_gnt,

  // Rx
  output  [C_DATA_WIDTH-1:0]                 m_axis_rx_tdata,
  output  [KEEP_WIDTH-1:0]                   m_axis_rx_tkeep,
  output                                     m_axis_rx_tlast,
  output                                     m_axis_rx_tvalid,
  input                                      m_axis_rx_tready,
  output  [21:0]                             m_axis_rx_tuser,
  input                                      rx_np_ok,
  input                                      rx_np_req,

  // Flow Control
  output  [11:0]                             fc_cpld,
  output  [7:0]                              fc_cplh,
  output  [11:0]                             fc_npd,
  output  [7:0]                              fc_nph,
  output  [11:0]                             fc_pd,
  output  [7:0]                              fc_ph,
  input   [2:0]                              fc_sel,

  input wire   [1:0]   pl_directed_link_change,
  input wire   [1:0]   pl_directed_link_width,
  input wire           pl_directed_link_speed,
  input wire           pl_directed_link_auton,
  input wire           pl_upstream_prefer_deemph,
  input wire           pl_downstream_deemph_source,
  input wire           pl_directed_ltssm_new_vld,
  input wire   [5:0]   pl_directed_ltssm_new,
  input wire           pl_directed_ltssm_stall,

  input wire           cm_rst_n,
  input wire           func_lvl_rst_n,
  input wire           pl_transmit_hot_rst,
  input wire   [31:0]  cfg_mgmt_di,
  input wire   [3:0]   cfg_mgmt_byte_en_n,
  input wire   [9:0]   cfg_mgmt_dwaddr,
  input wire           cfg_mgmt_wr_rw1c_as_rw_n,
  input wire           cfg_mgmt_wr_readonly_n,
  input wire           cfg_mgmt_wr_en_n,
  input wire           cfg_mgmt_rd_en_n,
  input wire           cfg_err_malformed_n,
  input wire           cfg_err_cor_n,
  input wire           cfg_err_ur_n,
  input wire           cfg_err_ecrc_n,
  input wire           cfg_err_cpl_timeout_n,
  input wire           cfg_err_cpl_abort_n,
  input wire           cfg_err_cpl_unexpect_n,
  input wire           cfg_err_poisoned_n,
  input wire           cfg_err_acs_n,
  input wire           cfg_err_atomic_egress_blocked_n,
  input wire           cfg_err_mc_blocked_n,
  input wire           cfg_err_internal_uncor_n,
  input wire           cfg_err_internal_cor_n,
  input wire           cfg_err_posted_n,
  input wire           cfg_err_locked_n,
  input wire           cfg_err_norecovery_n,
  input wire   [127:0] cfg_err_aer_headerlog,
  input wire   [47:0]  cfg_err_tlp_cpl_header,
  input wire           cfg_interrupt_n,
  input wire   [7:0]   cfg_interrupt_di,
  input wire           cfg_interrupt_assert_n,
  input wire           cfg_interrupt_stat_n,
  input wire   [7:0]   cfg_ds_bus_number,
  input wire   [4:0]   cfg_ds_device_number,
  input wire   [2:0]   cfg_ds_function_number,
  input wire   [7:0]   cfg_port_number,
  input wire           cfg_pm_halt_aspm_l0s_n,
  input wire           cfg_pm_halt_aspm_l1_n,
  input wire           cfg_pm_force_state_en_n,
  input wire   [1:0]   cfg_pm_force_state,
  input wire           cfg_pm_wake_n,
  input wire           cfg_turnoff_ok,
  input wire           cfg_pm_send_pme_to_n,
  input wire   [4:0]   cfg_pciecap_interrupt_msgnum,
  input wire           cfg_trn_pending,
  input wire   [2:0]   cfg_force_mps,
  input wire           cfg_force_common_clock_off,
  input wire           cfg_force_extended_sync_on,
  input wire   [63:0]  cfg_dsn,
  input wire   [4:0]   cfg_aer_interrupt_msgnum,
  input wire   [15:0]  cfg_dev_id,
  input wire   [15:0]  cfg_vend_id,
  input wire   [7:0]   cfg_rev_id,
  input wire   [15:0]  cfg_subsys_id,
  input wire   [15:0]  cfg_subsys_vend_id,
  input wire           drp_clk,
  input wire           drp_en,
  input wire           drp_we,
  input wire   [8:0]   drp_addr,
  input wire   [15:0]  drp_di,
  input wire   [1:0]   dbg_mode,
  input wire           dbg_sub_mode,
  input wire   [2:0]   pl_dbg_mode ,

  output wire          pl_sel_lnk_rate,
  output wire  [1:0]   pl_sel_lnk_width,
  output wire  [5:0]   pl_ltssm_state,
  output wire  [1:0]   pl_lane_reversal_mode,
  output wire          pl_phy_lnk_up,
  output wire  [2:0]   pl_tx_pm_state,
  output wire  [1:0]   pl_rx_pm_state,
  output wire          pl_link_upcfg_cap,
  output wire          pl_link_gen2_cap,
  output wire          pl_link_partner_gen2_supported,
  output wire  [2:0]   pl_initial_link_width,
  output wire          pl_directed_change_done,
  output wire          pl_received_hot_rst,
  output wire          lnk_clk_en,
  output wire  [31:0]  cfg_mgmt_do,
  output wire          cfg_mgmt_rd_wr_done,
  output wire          cfg_err_aer_headerlog_set,
  output wire          cfg_err_cpl_rdy,
  output wire          cfg_interrupt_rdy,
  output wire  [2:0]   cfg_interrupt_mmenable,
  output wire          cfg_interrupt_msienable,
  output wire  [7:0]   cfg_interrupt_do,
  output wire          cfg_interrupt_msixenable,
  output wire          cfg_interrupt_msixfm,
  output wire  [7:0]   cfg_bus_number,
  output wire  [4:0]   cfg_device_number,
  output wire  [2:0]   cfg_function_number,
  output wire  [15:0]  cfg_status,
  output wire  [15:0]  cfg_command,
  output wire  [15:0]  cfg_dstatus,
  output wire  [15:0]  cfg_dcommand,
  output wire  [15:0]  cfg_lstatus,
  output wire  [15:0]  cfg_lcommand,
  output wire  [15:0]  cfg_dcommand2,
  output wire          cfg_received_func_lvl_rst,
  output wire          cfg_msg_received,
  output wire  [15:0]  cfg_msg_data,
  output wire          cfg_msg_received_err_cor,
  output wire          cfg_msg_received_err_non_fatal,
  output wire          cfg_msg_received_err_fatal,
  output wire          cfg_msg_received_assert_int_a,
  output wire          cfg_msg_received_deassert_int_a,
  output wire          cfg_msg_received_assert_int_b,
  output wire          cfg_msg_received_deassert_int_b,
  output wire          cfg_msg_received_assert_int_c,
  output wire          cfg_msg_received_deassert_int_c,
  output wire          cfg_msg_received_assert_int_d,
  output wire          cfg_msg_received_deassert_int_d,
  output wire          cfg_msg_received_pm_pme,
  output wire          cfg_msg_received_pme_to_ack,
  output wire          cfg_msg_received_pme_to,
  output wire          cfg_msg_received_setslotpowerlimit,
  output wire          cfg_msg_received_unlock,
  output wire          cfg_msg_received_pm_as_nak,
  output wire          cfg_to_turnoff,
  output wire  [2:0]   cfg_pcie_link_state,
  output wire          cfg_pm_rcv_as_req_l1_n,
  output wire          cfg_pm_rcv_enter_l1_n,
  output wire          cfg_pm_rcv_enter_l23_n,
  output wire          cfg_pm_rcv_req_ack_n,
  output wire  [1:0]   cfg_pmcsr_powerstate,
  output wire          cfg_pmcsr_pme_en,
  output wire          cfg_pmcsr_pme_status,
  output wire          cfg_transaction,
  output wire          cfg_transaction_type,
  output wire  [6:0]   cfg_transaction_addr,
  output wire          cfg_command_io_enable,
  output wire          cfg_command_mem_enable,
  output wire          cfg_command_bus_master_enable,
  output wire          cfg_command_interrupt_disable,
  output wire          cfg_command_serr_en,
  output wire          cfg_bridge_serr_en,
  output wire          cfg_dev_status_corr_err_detected,
  output wire          cfg_dev_status_non_fatal_err_detected,
  output wire          cfg_dev_status_fatal_err_detected,
  output wire          cfg_dev_status_ur_detected,
  output wire          cfg_dev_control_corr_err_reporting_en,
  output wire          cfg_dev_control_non_fatal_reporting_en,
  output wire          cfg_dev_control_fatal_err_reporting_en,
  output wire          cfg_dev_control_ur_err_reporting_en,
  output wire          cfg_dev_control_enable_ro,
  output wire  [2:0]   cfg_dev_control_max_payload,
  output wire          cfg_dev_control_ext_tag_en,
  output wire          cfg_dev_control_phantom_en,
  output wire          cfg_dev_control_aux_power_en,
  output wire          cfg_dev_control_no_snoop_en,
  output wire  [2:0]   cfg_dev_control_max_read_req,
  output wire  [1:0]   cfg_link_status_current_speed,
  output wire  [3:0]   cfg_link_status_negotiated_width,
  output wire          cfg_link_status_link_training,
  output wire          cfg_link_status_dll_active,
  output wire          cfg_link_status_bandwidth_status,
  output wire          cfg_link_status_auto_bandwidth_status,
  output wire  [1:0]   cfg_link_control_aspm_control,
  output wire          cfg_link_control_rcb,
  output wire          cfg_link_control_link_disable,
  output wire          cfg_link_control_retrain_link,
  output wire          cfg_link_control_common_clock,
  output wire          cfg_link_control_extended_sync,
  output wire          cfg_link_control_clock_pm_en,
  output wire          cfg_link_control_hw_auto_width_dis,
  output wire          cfg_link_control_bandwidth_int_en,
  output wire          cfg_link_control_auto_bandwidth_int_en,
  output wire  [3:0]   cfg_dev_control2_cpl_timeout_val,
  output wire          cfg_dev_control2_cpl_timeout_dis,
  output wire          cfg_dev_control2_ari_forward_en,
  output wire          cfg_dev_control2_atomic_requester_en,
  output wire          cfg_dev_control2_atomic_egress_block,
  output wire          cfg_dev_control2_ido_req_en,
  output wire          cfg_dev_control2_ido_cpl_en,
  output wire          cfg_dev_control2_ltr_en,
  output wire          cfg_dev_control2_tlp_prefix_block,
  output wire          cfg_slot_control_electromech_il_ctl_pulse,
  output wire          cfg_root_control_syserr_corr_err_en,
  output wire          cfg_root_control_syserr_non_fatal_err_en,
  output wire          cfg_root_control_syserr_fatal_err_en,
  output wire          cfg_root_control_pme_int_en,
  output wire          cfg_aer_ecrc_check_en,
  output wire          cfg_aer_ecrc_gen_en,
  output wire          cfg_aer_rooterr_corr_err_reporting_en,
  output wire          cfg_aer_rooterr_non_fatal_err_reporting_en,
  output wire          cfg_aer_rooterr_fatal_err_reporting_en,
  output wire          cfg_aer_rooterr_corr_err_received,
  output wire          cfg_aer_rooterr_non_fatal_err_received,
  output wire          cfg_aer_rooterr_fatal_err_received,
  output wire  [6:0]   cfg_vc_tcvc_map,
  output wire          drp_rdy,
  output wire  [15:0]  drp_do,
  output wire  [63:0]  dbg_vec_a,
  output wire  [63:0]  dbg_vec_b,
  output wire  [11:0]  dbg_vec_c,
  output wire          dbg_sclr_a,
  output wire          dbg_sclr_b,
  output wire          dbg_sclr_c,
  output wire          dbg_sclr_d,
  output wire          dbg_sclr_e,
  output wire          dbg_sclr_f,
  output wire          dbg_sclr_g,
  output wire          dbg_sclr_h,
  output wire          dbg_sclr_i,
  output wire          dbg_sclr_j,
  output wire          dbg_sclr_k,
  output wire  [63:0]  trn_rdllp_data,
  output wire   [1:0]  trn_rdllp_src_rdy,
  output wire  [11:0]  pl_dbg_vec,

  input                       phy_rdy_n,
  input                       pipe_clk,
  input                       user_clk,
  input                       user_clk2,
  output wire                 pipe_rx0_polarity_gt,
  output wire                 pipe_rx1_polarity_gt,
  output wire                 pipe_rx2_polarity_gt,
  output wire                 pipe_rx3_polarity_gt,
  output wire                 pipe_rx4_polarity_gt,
  output wire                 pipe_rx5_polarity_gt,
  output wire                 pipe_rx6_polarity_gt,
  output wire                 pipe_rx7_polarity_gt,
  output wire                 pipe_tx_deemph_gt,
  output wire [2:0]           pipe_tx_margin_gt,
  output wire                 pipe_tx_rate_gt,
  output wire                 pipe_tx_rcvr_det_gt,
  output wire [1:0]           pipe_tx0_char_is_k_gt,
  output wire                 pipe_tx0_compliance_gt,
  output wire [15:0]          pipe_tx0_data_gt,
  output wire                 pipe_tx0_elec_idle_gt,
  output wire [1:0]           pipe_tx0_powerdown_gt,
  output wire [1:0]           pipe_tx1_char_is_k_gt,
  output wire                 pipe_tx1_compliance_gt,
  output wire [15:0]          pipe_tx1_data_gt,
  output wire                 pipe_tx1_elec_idle_gt,
  output wire [1:0]           pipe_tx1_powerdown_gt,
  output wire [1:0]           pipe_tx2_char_is_k_gt,
  output wire                 pipe_tx2_compliance_gt,
  output wire [15:0]          pipe_tx2_data_gt,
  output wire                 pipe_tx2_elec_idle_gt,
  output wire [1:0]           pipe_tx2_powerdown_gt,
  output wire [1:0]           pipe_tx3_char_is_k_gt,
  output wire                 pipe_tx3_compliance_gt,
  output wire [15:0]          pipe_tx3_data_gt,
  output wire                 pipe_tx3_elec_idle_gt,
  output wire [1:0]           pipe_tx3_powerdown_gt,
  output wire [1:0]           pipe_tx4_char_is_k_gt,
  output wire                 pipe_tx4_compliance_gt,
  output wire [15:0]          pipe_tx4_data_gt,
  output wire                 pipe_tx4_elec_idle_gt,
  output wire [1:0]           pipe_tx4_powerdown_gt,
  output wire [1:0]           pipe_tx5_char_is_k_gt,
  output wire                 pipe_tx5_compliance_gt,
  output wire [15:0]          pipe_tx5_data_gt,
  output wire                 pipe_tx5_elec_idle_gt,
  output wire [1:0]           pipe_tx5_powerdown_gt,
  output wire [1:0]           pipe_tx6_char_is_k_gt,
  output wire                 pipe_tx6_compliance_gt,
  output wire [15:0]          pipe_tx6_data_gt,
  output wire                 pipe_tx6_elec_idle_gt,
  output wire [1:0]           pipe_tx6_powerdown_gt,
  output wire [1:0]           pipe_tx7_char_is_k_gt,
  output wire                 pipe_tx7_compliance_gt,
  output wire [15:0]          pipe_tx7_data_gt,
  output wire                 pipe_tx7_elec_idle_gt,
  output wire [1:0]           pipe_tx7_powerdown_gt,

  input wire                 pipe_rx0_chanisaligned_gt,
  input wire  [1:0]          pipe_rx0_char_is_k_gt,
  input wire  [15:0]         pipe_rx0_data_gt,
  input wire                 pipe_rx0_elec_idle_gt,
  input wire                 pipe_rx0_phy_status_gt,
  input wire  [2:0]          pipe_rx0_status_gt,
  input wire                 pipe_rx0_valid_gt,
  input wire                 pipe_rx1_chanisaligned_gt,
  input wire  [1:0]          pipe_rx1_char_is_k_gt,
  input wire  [15:0]         pipe_rx1_data_gt,
  input wire                 pipe_rx1_elec_idle_gt,
  input wire                 pipe_rx1_phy_status_gt,
  input wire  [2:0]          pipe_rx1_status_gt,
  input wire                 pipe_rx1_valid_gt,
  input wire                 pipe_rx2_chanisaligned_gt,
  input wire  [1:0]          pipe_rx2_char_is_k_gt,
  input wire  [15:0]         pipe_rx2_data_gt,
  input wire                 pipe_rx2_elec_idle_gt,
  input wire                 pipe_rx2_phy_status_gt,
  input wire  [2:0]          pipe_rx2_status_gt,
  input wire                 pipe_rx2_valid_gt,
  input wire                 pipe_rx3_chanisaligned_gt,
  input wire  [1:0]          pipe_rx3_char_is_k_gt,
  input wire  [15:0]         pipe_rx3_data_gt,
  input wire                 pipe_rx3_elec_idle_gt,
  input wire                 pipe_rx3_phy_status_gt,
  input wire  [2:0]          pipe_rx3_status_gt,
  input wire                 pipe_rx3_valid_gt,
  input wire                 pipe_rx4_chanisaligned_gt,
  input wire  [1:0]          pipe_rx4_char_is_k_gt,
  input wire  [15:0]         pipe_rx4_data_gt,
  input wire                 pipe_rx4_elec_idle_gt,
  input wire                 pipe_rx4_phy_status_gt,
  input wire  [2:0]          pipe_rx4_status_gt,
  input wire                 pipe_rx4_valid_gt,
  input wire                 pipe_rx5_chanisaligned_gt,
  input wire  [1:0]          pipe_rx5_char_is_k_gt,
  input wire  [15:0]         pipe_rx5_data_gt,
  input wire                 pipe_rx5_elec_idle_gt,
  input wire                 pipe_rx5_phy_status_gt,
  input wire  [2:0]          pipe_rx5_status_gt,
  input wire                 pipe_rx5_valid_gt,
  input wire                 pipe_rx6_chanisaligned_gt,
  input wire  [1:0]          pipe_rx6_char_is_k_gt,
  input wire  [15:0]         pipe_rx6_data_gt,
  input wire                 pipe_rx6_elec_idle_gt,
  input wire                 pipe_rx6_phy_status_gt,
  input wire  [2:0]          pipe_rx6_status_gt,
  input wire                 pipe_rx6_valid_gt,
  input wire                 pipe_rx7_chanisaligned_gt,
  input wire  [1:0]          pipe_rx7_char_is_k_gt,
  input wire  [15:0]         pipe_rx7_data_gt,
  input wire                 pipe_rx7_elec_idle_gt,
  input wire                 pipe_rx7_phy_status_gt,
  input wire  [2:0]          pipe_rx7_status_gt,
  input wire                 pipe_rx7_valid_gt
);

  //wire declaration

  // TRN Interface
  wire [C_DATA_WIDTH-1:0]  trn_td;
  wire [REM_WIDTH-1:0]     trn_trem;
  wire                     trn_tsof;
  wire                     trn_teof;
  wire                     trn_tsrc_rdy;
  wire                     trn_tsrc_dsc;
  wire                     trn_terrfwd;
  wire                     trn_tecrc_gen;
  wire                     trn_tstr;
  wire                     trn_tcfg_gnt;
  wire                     trn_tdst_rdy;


  wire [127:0]  trn_rd;
  wire [1:0]     trn_rrem;
  wire                     trn_rdst_rdy;
  wire                     trn_rsof;
  wire                     trn_reof;
  wire                     trn_rsrc_rdy;
  wire                     trn_rsrc_dsc;
  wire                     trn_recrc_err;
  wire                     trn_rerrfwd;
  wire [7:0]               trn_rbar_hit;

  wire                 sys_reset_n_d;
  wire [1:0]           pipe_rx0_char_is_k;
  wire [1:0]           pipe_rx1_char_is_k;
  wire [1:0]           pipe_rx2_char_is_k;
  wire [1:0]           pipe_rx3_char_is_k;
  wire [1:0]           pipe_rx4_char_is_k;
  wire [1:0]           pipe_rx5_char_is_k;
  wire [1:0]           pipe_rx6_char_is_k;
  wire [1:0]           pipe_rx7_char_is_k;
  wire                 pipe_rx0_valid;
  wire                 pipe_rx1_valid;
  wire                 pipe_rx2_valid;
  wire                 pipe_rx3_valid;
  wire                 pipe_rx4_valid;
  wire                 pipe_rx5_valid;
  wire                 pipe_rx6_valid;
  wire                 pipe_rx7_valid;
  wire [15:0]          pipe_rx0_data;
  wire [15:0]          pipe_rx1_data;
  wire [15:0]          pipe_rx2_data;
  wire [15:0]          pipe_rx3_data;
  wire [15:0]          pipe_rx4_data;
  wire [15:0]          pipe_rx5_data;
  wire [15:0]          pipe_rx6_data;
  wire [15:0]          pipe_rx7_data;
  wire                 pipe_rx0_chanisaligned;
  wire                 pipe_rx1_chanisaligned;
  wire                 pipe_rx2_chanisaligned;
  wire                 pipe_rx3_chanisaligned;
  wire                 pipe_rx4_chanisaligned;
  wire                 pipe_rx5_chanisaligned;
  wire                 pipe_rx6_chanisaligned;
  wire                 pipe_rx7_chanisaligned;
  wire [2:0]           pipe_rx0_status;
  wire [2:0]           pipe_rx1_status;
  wire [2:0]           pipe_rx2_status;
  wire [2:0]           pipe_rx3_status;
  wire [2:0]           pipe_rx4_status;
  wire [2:0]           pipe_rx5_status;
  wire [2:0]           pipe_rx6_status;
  wire [2:0]           pipe_rx7_status;
  wire                 pipe_rx0_phy_status;
  wire                 pipe_rx1_phy_status;
  wire                 pipe_rx2_phy_status;
  wire                 pipe_rx3_phy_status;
  wire                 pipe_rx4_phy_status;
  wire                 pipe_rx5_phy_status;
  wire                 pipe_rx6_phy_status;
  wire                 pipe_rx7_phy_status;

  wire                 pipe_rx0_elec_idle;
  wire                 pipe_rx1_elec_idle;
  wire                 pipe_rx2_elec_idle;
  wire                 pipe_rx3_elec_idle;
  wire                 pipe_rx4_elec_idle;
  wire                 pipe_rx5_elec_idle;
  wire                 pipe_rx6_elec_idle;
  wire                 pipe_rx7_elec_idle;


  wire                 pipe_tx_reset;
  wire                 pipe_tx_rcvr_det;
  wire                 pipe_tx_rate;
  wire                 pipe_tx_deemph;
  wire [2:0]           pipe_tx_margin;
  wire                 pipe_rx0_polarity;
  wire                 pipe_rx1_polarity;
  wire                 pipe_rx2_polarity;
  wire                 pipe_rx3_polarity;
  wire                 pipe_rx4_polarity;
  wire                 pipe_rx5_polarity;
  wire                 pipe_rx6_polarity;
  wire                 pipe_rx7_polarity;
  wire                 pipe_tx0_compliance;
  wire                 pipe_tx1_compliance;
  wire                 pipe_tx2_compliance;
  wire                 pipe_tx3_compliance;
  wire                 pipe_tx4_compliance;
  wire                 pipe_tx5_compliance;
  wire                 pipe_tx6_compliance;
  wire                 pipe_tx7_compliance;
  wire [1:0]           pipe_tx0_char_is_k;
  wire [1:0]           pipe_tx1_char_is_k;
  wire [1:0]           pipe_tx2_char_is_k;
  wire [1:0]           pipe_tx3_char_is_k;
  wire [1:0]           pipe_tx4_char_is_k;
  wire [1:0]           pipe_tx5_char_is_k;
  wire [1:0]           pipe_tx6_char_is_k;
  wire [1:0]           pipe_tx7_char_is_k;
  wire [15:0]          pipe_tx0_data;
  wire [15:0]          pipe_tx1_data;
  wire [15:0]          pipe_tx2_data;
  wire [15:0]          pipe_tx3_data;
  wire [15:0]          pipe_tx4_data;
  wire [15:0]          pipe_tx5_data;
  wire [15:0]          pipe_tx6_data;
  wire [15:0]          pipe_tx7_data;
  wire                 pipe_tx0_elec_idle;
  wire                 pipe_tx1_elec_idle;
  wire                 pipe_tx2_elec_idle;
  wire                 pipe_tx3_elec_idle;
  wire                 pipe_tx4_elec_idle;
  wire                 pipe_tx5_elec_idle;
  wire                 pipe_tx6_elec_idle;
  wire                 pipe_tx7_elec_idle;
  wire [1:0]           pipe_tx0_powerdown;
  wire [1:0]           pipe_tx1_powerdown;
  wire [1:0]           pipe_tx2_powerdown;
  wire [1:0]           pipe_tx3_powerdown;
  wire [1:0]           pipe_tx4_powerdown;
  wire [1:0]           pipe_tx5_powerdown;
  wire [1:0]           pipe_tx6_powerdown;
  wire [1:0]           pipe_tx7_powerdown;

  wire                 cfg_received_func_lvl_rst_n;
  wire                 cfg_err_cpl_rdy_n;
  wire                 cfg_interrupt_rdy_n;
  reg [7:0]            cfg_bus_number_d;
  reg [4:0]            cfg_device_number_d;
  reg [2:0]            cfg_function_number_d;

  wire                 cfg_mgmt_rd_wr_done_n;
  wire                 pl_phy_lnk_up_n;
  wire                 cfg_err_aer_headerlog_set_n;
  wire                 cfg_turnoff_ok_w;

  assign        cfg_received_func_lvl_rst = ~cfg_received_func_lvl_rst_n;

  assign        cfg_err_cpl_rdy = ~cfg_err_cpl_rdy_n;

  assign        cfg_interrupt_rdy = ~cfg_interrupt_rdy_n;

  assign        cfg_mgmt_rd_wr_done = ~cfg_mgmt_rd_wr_done_n;

  assign        pl_phy_lnk_up = ~pl_phy_lnk_up_n;

  assign        cfg_err_aer_headerlog_set = ~cfg_err_aer_headerlog_set_n;

  assign        cfg_to_turnoff = cfg_msg_received_pme_to;

  assign        cfg_status   = {16'b0};

  assign        cfg_command  = {5'b0,
                                cfg_command_interrupt_disable,
                                1'b0,
                                cfg_command_serr_en,
                                5'b0,
                                cfg_command_bus_master_enable,
                                cfg_command_mem_enable,
                                cfg_command_io_enable};

  assign        cfg_dstatus  = {10'h0,
                                cfg_trn_pending,
                                1'b0,
                                cfg_dev_status_ur_detected,
                                cfg_dev_status_fatal_err_detected,
                                cfg_dev_status_non_fatal_err_detected,
                                cfg_dev_status_corr_err_detected};

  assign        cfg_dcommand = {1'b0,
                                cfg_dev_control_max_read_req,
                                cfg_dev_control_no_snoop_en,
                                cfg_dev_control_aux_power_en,
                                cfg_dev_control_phantom_en,
                                cfg_dev_control_ext_tag_en,
                                cfg_dev_control_max_payload,
                                cfg_dev_control_enable_ro,
                                cfg_dev_control_ur_err_reporting_en,
                                cfg_dev_control_fatal_err_reporting_en,
                                cfg_dev_control_non_fatal_reporting_en,
                                cfg_dev_control_corr_err_reporting_en };

  assign        cfg_lstatus  = {cfg_link_status_auto_bandwidth_status,
                                cfg_link_status_bandwidth_status,
                                cfg_link_status_dll_active,
                                (LINK_STATUS_SLOT_CLOCK_CONFIG == "TRUE") ? 1'b1 : 1'b0,
                                cfg_link_status_link_training,
                                1'b0,
                                {2'b00, cfg_link_status_negotiated_width},
                                {2'b00, cfg_link_status_current_speed} };

  assign        cfg_lcommand = {4'b0,
                                cfg_link_control_auto_bandwidth_int_en,
                                cfg_link_control_bandwidth_int_en,
                                cfg_link_control_hw_auto_width_dis,
                                cfg_link_control_clock_pm_en,
                                cfg_link_control_extended_sync,
                                cfg_link_control_common_clock,
                                cfg_link_control_retrain_link,
                                cfg_link_control_link_disable,
                                cfg_link_control_rcb,
                                1'b0,
                                cfg_link_control_aspm_control};

  assign       cfg_bus_number = cfg_bus_number_d;

  assign       cfg_device_number = cfg_device_number_d;

  assign       cfg_function_number =  cfg_function_number_d;

  assign       cfg_dcommand2 = {4'b0,
                                cfg_dev_control2_tlp_prefix_block,
                                cfg_dev_control2_ltr_en,
                                cfg_dev_control2_ido_cpl_en,
                                cfg_dev_control2_ido_req_en,
                                cfg_dev_control2_atomic_egress_block,
                                cfg_dev_control2_atomic_requester_en,
                                cfg_dev_control2_ari_forward_en,
                                cfg_dev_control2_cpl_timeout_dis,
                                cfg_dev_control2_cpl_timeout_val};

  // Capture Bus/Device/Function number

  always @(posedge user_clk_out) begin
    if (~user_lnk_up)
    begin
      cfg_bus_number_d <= 8'b0;
    end // if (~user_lnk_up)
    else if (~cfg_msg_received)
    begin
      cfg_bus_number_d <= cfg_msg_data[15:8];
    end // if (~cfg_msg_received)
  end

  always @(posedge user_clk_out) begin
    if (~user_lnk_up)
    begin
      cfg_device_number_d <= 5'b0;
    end // if (~user_lnk_up)
    else if (~cfg_msg_received)
    begin
      cfg_device_number_d <= cfg_msg_data[7:3];
    end // if (~cfg_msg_received)
  end

  always @(posedge user_clk_out) begin
    if (~user_lnk_up)
    begin
      cfg_function_number_d <= 3'b0;
    end // if (~user_lnk_up)
    else if (~cfg_msg_received)
    begin
      cfg_function_number_d <= cfg_msg_data[2:0];
    end // if (~cfg_msg_received)
  end

model_ap2_tst_axi_basic_top #(
  .C_DATA_WIDTH     (C_DATA_WIDTH),       // RX/TX interface data width
  .C_FAMILY         ("X7"),               // Targeted FPGA family
  .C_ROOT_PORT      ("FALSE"),            // PCIe block is in root port mode
  .C_PM_PRIORITY    ("FALSE")             // Disable TX packet boundary thrtl

  ) model_ap2_tst_axi_basic_top (
    //---------------------------------------------//
    // User Design I/O                             //
    //---------------------------------------------//

    // AXI TX
    //-----------
    .s_axis_tx_tdata          (s_axis_tx_tdata),          //  input
    .s_axis_tx_tvalid         (s_axis_tx_tvalid),         //  input
    .s_axis_tx_tready         (s_axis_tx_tready),         //  output
    .s_axis_tx_tkeep          (s_axis_tx_tkeep),          //  input
    .s_axis_tx_tlast          (s_axis_tx_tlast),          //  input
    .s_axis_tx_tuser          (s_axis_tx_tuser),          //  input

    // AXI RX
    //-----------
    .m_axis_rx_tdata          (m_axis_rx_tdata),          //  output
    .m_axis_rx_tvalid         (m_axis_rx_tvalid),         //  output
    .m_axis_rx_tready         (m_axis_rx_tready),         //  input
    .m_axis_rx_tkeep          (m_axis_rx_tkeep),          //  output
    .m_axis_rx_tlast          (m_axis_rx_tlast),          //  output
    .m_axis_rx_tuser          (m_axis_rx_tuser),          //  output

    // User Misc.
    //-----------
    .user_turnoff_ok          (cfg_turnoff_ok),           //  input
    .user_tcfg_gnt            (tx_cfg_gnt),               //  input

    //---------------------------------------------//
    // PCIe Block I/O                              //
    //---------------------------------------------//

    // TRN TX
    //-----------
    .trn_td                   (trn_td),                   //  output
    .trn_tsof                 (trn_tsof),                 //  output
    .trn_teof                 (trn_teof),                 //  output
    .trn_tsrc_rdy             (trn_tsrc_rdy),             //  output
    .trn_tdst_rdy             (trn_tdst_rdy),             //  input
    .trn_tsrc_dsc             (trn_tsrc_dsc),             //  output
    .trn_trem                 (trn_trem),                 //  output
    .trn_terrfwd              (trn_terrfwd),              //  output
    .trn_tstr                 (trn_tstr),                 //  output
    .trn_tbuf_av              (tx_buf_av),                //  input
    .trn_tecrc_gen            (trn_tecrc_gen),            //  output

    // TRN RX
    //-----------
    .trn_rd                   (trn_rd),                   //  input
    .trn_rsof                 (trn_rsof),                 //  input
    .trn_reof                 (trn_reof),                 //  input
    .trn_rsrc_rdy             (trn_rsrc_rdy),             //  input
    .trn_rdst_rdy             (trn_rdst_rdy),             //  output
    .trn_rsrc_dsc             (trn_rsrc_dsc),             //  input
    .trn_rrem                 (trn_rrem),                 //  input
    .trn_rerrfwd              (trn_rerrfwd),              //  input
    .trn_rbar_hit             (trn_rbar_hit[6:0]),             //  input
    .trn_recrc_err            (trn_recrc_err),            //  input

    // TRN Misc.
    //-----------
    .trn_tcfg_req             ( tx_cfg_req ),             //  input
    .trn_tcfg_gnt             ( trn_tcfg_gnt),            //  output
    .trn_lnk_up               ( user_lnk_up),             //  input

    // Fuji3/Virtex6 PM
    //-----------
    .cfg_pcie_link_state      (cfg_pcie_link_state),      //  input

    // Virtex6 PM
    //-----------
    .cfg_pm_send_pme_to       (1'b0),                     //  input  NOT USED FOR EP
    .cfg_pmcsr_powerstate     (cfg_pmcsr_powerstate),     //  input
    .trn_rdllp_data           (32'b0),                    //  input - Not used in 7-series
    .trn_rdllp_src_rdy        (1'b0),                     //  input -- Not used in 7-series

    // Power Mgmt for S6/V6
    //-----------
    .cfg_to_turnoff           (cfg_to_turnoff),           //  input
    .cfg_turnoff_ok           (cfg_turnoff_ok_w),         //  output

    // System
    //-----------
    .user_clk                 (user_clk_out),             //  input
    .user_rst                 (user_reset),               //  input
    .np_counter               ()                          //  output

  );


 //-------------------------------------------------------
 // PCI Express Pipe Wrapper
 //-------------------------------------------------------
model_ap2_tst_pcie_7x # (
    .AER_BASE_PTR    ( AER_BASE_PTR ),
    .AER_CAP_ECRC_CHECK_CAPABLE      ( AER_CAP_ECRC_CHECK_CAPABLE ),
    .AER_CAP_ECRC_GEN_CAPABLE( AER_CAP_ECRC_GEN_CAPABLE ),
    .AER_CAP_ID      ( AER_CAP_ID ),
    .AER_CAP_MULTIHEADER ( AER_CAP_MULTIHEADER ),
    .AER_CAP_NEXTPTR ( AER_CAP_NEXTPTR ),
    .AER_CAP_ON      ( AER_CAP_ON ),
    .AER_CAP_OPTIONAL_ERR_SUPPORT    ( AER_CAP_OPTIONAL_ERR_SUPPORT ),
    .AER_CAP_PERMIT_ROOTERR_UPDATE   ( AER_CAP_PERMIT_ROOTERR_UPDATE ),
    .AER_CAP_VERSION ( AER_CAP_VERSION ),
    .ALLOW_X8_GEN2 (ALLOW_X8_GEN2),
    .BAR0    ( BAR0 ),
    .BAR1    ( BAR1 ),
    .BAR2    ( BAR2 ),
    .BAR3    ( BAR3 ),
    .BAR4    ( BAR4 ),
    .BAR5    ( BAR5 ),
    .C_DATA_WIDTH ( C_DATA_WIDTH ),
    .CAPABILITIES_PTR( CAPABILITIES_PTR ),
    .CFG_ECRC_ERR_CPLSTAT    ( CFG_ECRC_ERR_CPLSTAT ),
    .CARDBUS_CIS_POINTER     ( CARDBUS_CIS_POINTER ),
    .CLASS_CODE      ( CLASS_CODE ),
    .CMD_INTX_IMPLEMENTED    ( CMD_INTX_IMPLEMENTED ),
    .CPL_TIMEOUT_DISABLE_SUPPORTED   ( CPL_TIMEOUT_DISABLE_SUPPORTED ),
    .CPL_TIMEOUT_RANGES_SUPPORTED    ( CPL_TIMEOUT_RANGES_SUPPORTED ),
    .CRM_MODULE_RSTS (CRM_MODULE_RSTS),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE     ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE     ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE ),
    .DEV_CAP_ENDPOINT_L0S_LATENCY    ( DEV_CAP_ENDPOINT_L0S_LATENCY ),
    .DEV_CAP_ENDPOINT_L1_LATENCY     ( DEV_CAP_ENDPOINT_L1_LATENCY ),
    .DEV_CAP_EXT_TAG_SUPPORTED ( DEV_CAP_EXT_TAG_SUPPORTED ),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE    ( DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE ),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED   ( DEV_CAP_MAX_PAYLOAD_SUPPORTED ),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT ( DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT ),
    .DEV_CAP_ROLE_BASED_ERROR( DEV_CAP_ROLE_BASED_ERROR ),
    .DEV_CAP_RSVD_14_12      ( DEV_CAP_RSVD_14_12 ),
    .DEV_CAP_RSVD_17_16      ( DEV_CAP_RSVD_17_16 ),
    .DEV_CAP_RSVD_31_29      ( DEV_CAP_RSVD_31_29 ),
    .DEV_CONTROL_AUX_POWER_SUPPORTED ( DEV_CONTROL_AUX_POWER_SUPPORTED ),
    .DEV_CONTROL_EXT_TAG_DEFAULT ( DEV_CONTROL_EXT_TAG_DEFAULT ),
    .DISABLE_ASPM_L1_TIMER   ( DISABLE_ASPM_L1_TIMER ),
    .DISABLE_BAR_FILTERING   ( DISABLE_BAR_FILTERING ),
    .DISABLE_ID_CHECK( DISABLE_ID_CHECK ),
    .DISABLE_LANE_REVERSAL   ( DISABLE_LANE_REVERSAL ),
    .DISABLE_RX_POISONED_RESP (DISABLE_RX_POISONED_RESP),
    .DISABLE_RX_TC_FILTER    ( DISABLE_RX_TC_FILTER ),
    .DISABLE_SCRAMBLING      ( DISABLE_SCRAMBLING ),
    .DNSTREAM_LINK_NUM ( DNSTREAM_LINK_NUM ),
    .DSN_BASE_PTR    ( DSN_BASE_PTR ),
    .DSN_CAP_ID      ( DSN_CAP_ID ),
    .DSN_CAP_NEXTPTR ( DSN_CAP_NEXTPTR ),
    .DSN_CAP_ON      ( DSN_CAP_ON ),
    .DSN_CAP_VERSION ( DSN_CAP_VERSION ),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED(DEV_CAP2_ARI_FORWARDING_SUPPORTED),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED (DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED (DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED (DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED (DEV_CAP2_CAS128_COMPLETER_SUPPORTED),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED (DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED (DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED (DEV_CAP2_LTR_MECHANISM_SUPPORTED),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES (DEV_CAP2_MAX_ENDEND_TLP_PREFIXES),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING (DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED (DEV_CAP2_TPH_COMPLETER_SUPPORTED),
    .DISABLE_ERR_MSG (DISABLE_ERR_MSG),
    .DISABLE_LOCKED_FILTER (DISABLE_LOCKED_FILTER),
    .DISABLE_PPM_FILTER (DISABLE_PPM_FILTER),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED (ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED),
    .ENABLE_MSG_ROUTE( ENABLE_MSG_ROUTE ),
    .ENABLE_RX_TD_ECRC_TRIM  ( ENABLE_RX_TD_ECRC_TRIM ),
    .ENTER_RVRY_EI_L0( ENTER_RVRY_EI_L0 ),
    .EXIT_LOOPBACK_ON_EI (EXIT_LOOPBACK_ON_EI),
    .EXPANSION_ROM   ( EXPANSION_ROM ),
    .EXT_CFG_CAP_PTR ( EXT_CFG_CAP_PTR ),
    .EXT_CFG_XP_CAP_PTR      ( EXT_CFG_XP_CAP_PTR ),
    .HEADER_TYPE     ( HEADER_TYPE ),
    .INFER_EI( INFER_EI ),
    .INTERRUPT_PIN   ( INTERRUPT_PIN ),
    .INTERRUPT_STAT_AUTO (INTERRUPT_STAT_AUTO),
    .IS_SWITCH ( IS_SWITCH ),
    .LAST_CONFIG_DWORD ( LAST_CONFIG_DWORD ),
    .LINK_CAP_ASPM_OPTIONALITY ( LINK_CAP_ASPM_OPTIONALITY ),
    .LINK_CAP_ASPM_SUPPORT   ( LINK_CAP_ASPM_SUPPORT ),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT ( LINK_CAP_CLOCK_POWER_MANAGEMENT ),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP  ( LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1   ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2   ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1  ( LINK_CAP_L0S_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2  ( LINK_CAP_L0S_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1    ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2    ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1   ( LINK_CAP_L1_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2   ( LINK_CAP_L1_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP (LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP),
    .LINK_CAP_MAX_LINK_SPEED ( LINK_CAP_MAX_LINK_SPEED ),
    .LINK_CAP_MAX_LINK_WIDTH ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_RSVD_23( LINK_CAP_RSVD_23 ),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE    ( LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE ),
    .LINK_CONTROL_RCB( LINK_CONTROL_RCB ),
    .LINK_CTRL2_DEEMPHASIS   ( LINK_CTRL2_DEEMPHASIS ),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE  ( LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE ),
    .LINK_CTRL2_TARGET_LINK_SPEED    ( LINK_CTRL2_TARGET_LINK_SPEED ),
    .LINK_STATUS_SLOT_CLOCK_CONFIG   ( LINK_STATUS_SLOT_CLOCK_CONFIG ),
    .LL_ACK_TIMEOUT  ( LL_ACK_TIMEOUT ),
    .LL_ACK_TIMEOUT_EN ( LL_ACK_TIMEOUT_EN ),
    .LL_ACK_TIMEOUT_FUNC     ( LL_ACK_TIMEOUT_FUNC ),
    .LL_REPLAY_TIMEOUT ( LL_REPLAY_TIMEOUT ),
    .LL_REPLAY_TIMEOUT_EN    ( LL_REPLAY_TIMEOUT_EN ),
    .LL_REPLAY_TIMEOUT_FUNC  ( LL_REPLAY_TIMEOUT_FUNC ),
    .LTSSM_MAX_LINK_WIDTH    ( LTSSM_MAX_LINK_WIDTH ),
    .MPS_FORCE (MPS_FORCE),
    .MSI_BASE_PTR    ( MSI_BASE_PTR ),
    .MSI_CAP_ID      ( MSI_CAP_ID ),
    .MSI_CAP_MULTIMSGCAP     ( MSI_CAP_MULTIMSGCAP ),
    .MSI_CAP_MULTIMSG_EXTENSION      ( MSI_CAP_MULTIMSG_EXTENSION ),
    .MSI_CAP_NEXTPTR ( MSI_CAP_NEXTPTR ),
    .MSI_CAP_ON      ( MSI_CAP_ON ),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE      ( MSI_CAP_PER_VECTOR_MASKING_CAPABLE ),
    .MSI_CAP_64_BIT_ADDR_CAPABLE     ( MSI_CAP_64_BIT_ADDR_CAPABLE ),
    .MSIX_BASE_PTR   ( MSIX_BASE_PTR ),
    .MSIX_CAP_ID     ( MSIX_CAP_ID ),
    .MSIX_CAP_NEXTPTR( MSIX_CAP_NEXTPTR ),
    .MSIX_CAP_ON     ( MSIX_CAP_ON ),
    .MSIX_CAP_PBA_BIR( MSIX_CAP_PBA_BIR ),
    .MSIX_CAP_PBA_OFFSET     ( MSIX_CAP_PBA_OFFSET ),
    .MSIX_CAP_TABLE_BIR      ( MSIX_CAP_TABLE_BIR ),
    .MSIX_CAP_TABLE_OFFSET   ( MSIX_CAP_TABLE_OFFSET ),
    .MSIX_CAP_TABLE_SIZE     ( MSIX_CAP_TABLE_SIZE ),
    .N_FTS_COMCLK_GEN1 ( N_FTS_COMCLK_GEN1 ),
    .N_FTS_COMCLK_GEN2 ( N_FTS_COMCLK_GEN2 ),
    .N_FTS_GEN1      ( N_FTS_GEN1 ),
    .N_FTS_GEN2      ( N_FTS_GEN2 ),
    .PCIE_BASE_PTR   ( PCIE_BASE_PTR ),
    .PCIE_CAP_CAPABILITY_ID  ( PCIE_CAP_CAPABILITY_ID ),
    .PCIE_CAP_CAPABILITY_VERSION     ( PCIE_CAP_CAPABILITY_VERSION ),
    .PCIE_CAP_DEVICE_PORT_TYPE ( PCIE_CAP_DEVICE_PORT_TYPE ),
    .PCIE_CAP_NEXTPTR( PCIE_CAP_NEXTPTR ),
    .PCIE_CAP_ON     ( PCIE_CAP_ON ),
    .PCIE_CAP_RSVD_15_14     ( PCIE_CAP_RSVD_15_14 ),
    .PCIE_CAP_SLOT_IMPLEMENTED ( PCIE_CAP_SLOT_IMPLEMENTED ),
    .PCIE_REVISION   ( PCIE_REVISION ),
    .PL_AUTO_CONFIG  ( PL_AUTO_CONFIG ),
    .PL_FAST_TRAIN   ( PL_FAST_TRAIN ),
    .PM_ASPML0S_TIMEOUT ( PM_ASPML0S_TIMEOUT ),
    .PM_ASPML0S_TIMEOUT_EN ( PM_ASPML0S_TIMEOUT_EN ),
    .PM_ASPML0S_TIMEOUT_FUNC ( PM_ASPML0S_TIMEOUT_FUNC ),
    .PM_ASPM_FASTEXIT ( PM_ASPM_FASTEXIT ),
    .PM_BASE_PTR     ( PM_BASE_PTR ),
    .PM_CAP_AUXCURRENT ( PM_CAP_AUXCURRENT ),
    .PM_CAP_D1SUPPORT( PM_CAP_D1SUPPORT ),
    .PM_CAP_D2SUPPORT( PM_CAP_D2SUPPORT ),
    .PM_CAP_DSI      ( PM_CAP_DSI ),
    .PM_CAP_ID ( PM_CAP_ID ),
    .PM_CAP_NEXTPTR  ( PM_CAP_NEXTPTR ),
    .PM_CAP_ON ( PM_CAP_ON ),
    .PM_CAP_PME_CLOCK( PM_CAP_PME_CLOCK ),
    .PM_CAP_PMESUPPORT ( PM_CAP_PMESUPPORT ),
    .PM_CAP_RSVD_04  ( PM_CAP_RSVD_04 ),
    .PM_CAP_VERSION  ( PM_CAP_VERSION ),
    .PM_CSR_B2B3     ( PM_CSR_B2B3 ),
    .PM_CSR_BPCCEN   ( PM_CSR_BPCCEN ),
    .PM_CSR_NOSOFTRST( PM_CSR_NOSOFTRST ),
    .PM_DATA0( PM_DATA0 ),
    .PM_DATA1( PM_DATA1 ),
    .PM_DATA2( PM_DATA2 ),
    .PM_DATA3( PM_DATA3 ),
    .PM_DATA4( PM_DATA4 ),
    .PM_DATA5( PM_DATA5 ),
    .PM_DATA6( PM_DATA6 ),
    .PM_DATA7( PM_DATA7 ),
    .PM_DATA_SCALE0  ( PM_DATA_SCALE0 ),
    .PM_DATA_SCALE1  ( PM_DATA_SCALE1 ),
    .PM_DATA_SCALE2  ( PM_DATA_SCALE2 ),
    .PM_DATA_SCALE3  ( PM_DATA_SCALE3 ),
    .PM_DATA_SCALE4  ( PM_DATA_SCALE4 ),
    .PM_DATA_SCALE5  ( PM_DATA_SCALE5 ),
    .PM_DATA_SCALE6  ( PM_DATA_SCALE6 ),
    .PM_DATA_SCALE7  ( PM_DATA_SCALE7 ),
    .PM_MF (PM_MF),
    .RBAR_BASE_PTR (RBAR_BASE_PTR),
    .RBAR_CAP_CONTROL_ENCODEDBAR0 (RBAR_CAP_CONTROL_ENCODEDBAR0),
    .RBAR_CAP_CONTROL_ENCODEDBAR1 (RBAR_CAP_CONTROL_ENCODEDBAR1),
    .RBAR_CAP_CONTROL_ENCODEDBAR2 (RBAR_CAP_CONTROL_ENCODEDBAR2),
    .RBAR_CAP_CONTROL_ENCODEDBAR3 (RBAR_CAP_CONTROL_ENCODEDBAR3),
    .RBAR_CAP_CONTROL_ENCODEDBAR4 (RBAR_CAP_CONTROL_ENCODEDBAR4),
    .RBAR_CAP_CONTROL_ENCODEDBAR5 (RBAR_CAP_CONTROL_ENCODEDBAR5),
    .RBAR_CAP_ID (RBAR_CAP_ID),
    .RBAR_CAP_INDEX0 (RBAR_CAP_INDEX0),
    .RBAR_CAP_INDEX1 (RBAR_CAP_INDEX1),
    .RBAR_CAP_INDEX2 (RBAR_CAP_INDEX2),
    .RBAR_CAP_INDEX3 (RBAR_CAP_INDEX3),
    .RBAR_CAP_INDEX4 (RBAR_CAP_INDEX4),
    .RBAR_CAP_INDEX5 (RBAR_CAP_INDEX5),
    .RBAR_CAP_NEXTPTR (RBAR_CAP_NEXTPTR),
    .RBAR_CAP_ON (RBAR_CAP_ON),
    .RBAR_CAP_SUP0 (RBAR_CAP_SUP0),
    .RBAR_CAP_SUP1 (RBAR_CAP_SUP1),
    .RBAR_CAP_SUP2 (RBAR_CAP_SUP2),
    .RBAR_CAP_SUP3 (RBAR_CAP_SUP3),
    .RBAR_CAP_SUP4 (RBAR_CAP_SUP4),
    .RBAR_CAP_SUP5 (RBAR_CAP_SUP5),
    .RBAR_CAP_VERSION (RBAR_CAP_VERSION),
    .RBAR_NUM (RBAR_NUM),
    .RECRC_CHK  (RECRC_CHK),
    .RECRC_CHK_TRIM (RECRC_CHK_TRIM),
    .ROOT_CAP_CRS_SW_VISIBILITY      ( ROOT_CAP_CRS_SW_VISIBILITY ),
    .RP_AUTO_SPD       ( RP_AUTO_SPD ),
    .RP_AUTO_SPD_LOOPCNT        ( RP_AUTO_SPD_LOOPCNT ),
    .SELECT_DLL_IF   ( SELECT_DLL_IF ),
    .SLOT_CAP_ATT_BUTTON_PRESENT     ( SLOT_CAP_ATT_BUTTON_PRESENT ),
    .SLOT_CAP_ATT_INDICATOR_PRESENT  ( SLOT_CAP_ATT_INDICATOR_PRESENT ),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT ( SLOT_CAP_ELEC_INTERLOCK_PRESENT ),
    .SLOT_CAP_HOTPLUG_CAPABLE( SLOT_CAP_HOTPLUG_CAPABLE ),
    .SLOT_CAP_HOTPLUG_SURPRISE ( SLOT_CAP_HOTPLUG_SURPRISE ),
    .SLOT_CAP_MRL_SENSOR_PRESENT     ( SLOT_CAP_MRL_SENSOR_PRESENT ),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT ( SLOT_CAP_NO_CMD_COMPLETED_SUPPORT ),
    .SLOT_CAP_PHYSICAL_SLOT_NUM      ( SLOT_CAP_PHYSICAL_SLOT_NUM ),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT ( SLOT_CAP_POWER_CONTROLLER_PRESENT ),
    .SLOT_CAP_POWER_INDICATOR_PRESENT( SLOT_CAP_POWER_INDICATOR_PRESENT ),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE ( SLOT_CAP_SLOT_POWER_LIMIT_SCALE ),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE ( SLOT_CAP_SLOT_POWER_LIMIT_VALUE ),
    .SPARE_BIT0      ( SPARE_BIT0 ),
    .SPARE_BIT1      ( SPARE_BIT1 ),
    .SPARE_BIT2      ( SPARE_BIT2 ),
    .SPARE_BIT3      ( SPARE_BIT3 ),
    .SPARE_BIT4      ( SPARE_BIT4 ),
    .SPARE_BIT5      ( SPARE_BIT5 ),
    .SPARE_BIT6      ( SPARE_BIT6 ),
    .SPARE_BIT7      ( SPARE_BIT7 ),
    .SPARE_BIT8      ( SPARE_BIT8 ),
    .SPARE_BYTE0     ( SPARE_BYTE0 ),
    .SPARE_BYTE1     ( SPARE_BYTE1 ),
    .SPARE_BYTE2     ( SPARE_BYTE2 ),
    .SPARE_BYTE3     ( SPARE_BYTE3 ),
    .SPARE_WORD0     ( SPARE_WORD0 ),
    .SPARE_WORD1     ( SPARE_WORD1 ),
    .SPARE_WORD2     ( SPARE_WORD2 ),
    .SPARE_WORD3     ( SPARE_WORD3 ),
    .SSL_MESSAGE_AUTO (SSL_MESSAGE_AUTO),
    .TECRC_EP_INV      ( TECRC_EP_INV ),
    .TL_RBYPASS(TL_RBYPASS),
    .TL_RX_RAM_RADDR_LATENCY ( TL_RX_RAM_RADDR_LATENCY ),
    .TL_RX_RAM_RDATA_LATENCY ( TL_RX_RAM_RDATA_LATENCY ),
    .TL_RX_RAM_WRITE_LATENCY ( TL_RX_RAM_WRITE_LATENCY ),
    .TL_TFC_DISABLE  ( TL_TFC_DISABLE ),
    .TL_TX_CHECKS_DISABLE    ( TL_TX_CHECKS_DISABLE ),
    .TL_TX_RAM_RADDR_LATENCY ( TL_TX_RAM_RADDR_LATENCY ),
    .TL_TX_RAM_RDATA_LATENCY ( TL_TX_RAM_RDATA_LATENCY ),
    .TL_TX_RAM_WRITE_LATENCY ( TL_TX_RAM_WRITE_LATENCY ),
    .TRN_DW (TRN_DW),
    .TRN_NP_FC (TRN_NP_FC),
    .UPCONFIG_CAPABLE( UPCONFIG_CAPABLE ),
    .UPSTREAM_FACING ( UPSTREAM_FACING ),
    .UR_ATOMIC (UR_ATOMIC),
    .UR_CFG1 (UR_CFG1),
    .UR_INV_REQ(UR_INV_REQ),
    .UR_PRS_RESPONSE (UR_PRS_RESPONSE),
    .USER_CLK2_DIV2 (USER_CLK2_DIV2),
    .USER_CLK_FREQ   ( USER_CLK_FREQ ),
    .USE_RID_PINS (USE_RID_PINS),
    .VC0_CPL_INFINITE( VC0_CPL_INFINITE ),
    .VC0_RX_RAM_LIMIT( VC0_RX_RAM_LIMIT ),
    .VC0_TOTAL_CREDITS_CD    ( VC0_TOTAL_CREDITS_CD ),
    .VC0_TOTAL_CREDITS_CH    ( VC0_TOTAL_CREDITS_CH ),
    .VC0_TOTAL_CREDITS_NPD (VC0_TOTAL_CREDITS_NPD),
    .VC0_TOTAL_CREDITS_NPH   ( VC0_TOTAL_CREDITS_NPH ),
    .VC0_TOTAL_CREDITS_PD    ( VC0_TOTAL_CREDITS_PD ),
    .VC0_TOTAL_CREDITS_PH    ( VC0_TOTAL_CREDITS_PH ),
    .VC0_TX_LASTPACKET ( VC0_TX_LASTPACKET ),
    .VC_BASE_PTR     ( VC_BASE_PTR ),
    .VC_CAP_ID ( VC_CAP_ID ),
    .VC_CAP_NEXTPTR  ( VC_CAP_NEXTPTR ),
    .VC_CAP_ON ( VC_CAP_ON ),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS( VC_CAP_REJECT_SNOOP_TRANSACTIONS ),
    .VC_CAP_VERSION  ( VC_CAP_VERSION ),
    .VSEC_BASE_PTR   ( VSEC_BASE_PTR ),
    .VSEC_CAP_HDR_ID ( VSEC_CAP_HDR_ID ),
    .VSEC_CAP_HDR_LENGTH     ( VSEC_CAP_HDR_LENGTH ),
    .VSEC_CAP_HDR_REVISION   ( VSEC_CAP_HDR_REVISION ),
    .VSEC_CAP_ID     ( VSEC_CAP_ID ),
    .VSEC_CAP_IS_LINK_VISIBLE( VSEC_CAP_IS_LINK_VISIBLE ),
    .VSEC_CAP_NEXTPTR( VSEC_CAP_NEXTPTR ),
    .VSEC_CAP_ON     ( VSEC_CAP_ON ),
    .VSEC_CAP_VERSION( VSEC_CAP_VERSION )
  ) model_ap2_tst_pcie_7x_i (
    .trn_lnk_up                                ( trn_lnk_up ),
    .trn_clk                                   ( user_clk_out ),
    .lnk_clk_en                                ( lnk_clk_en),
    .user_rst_n                                ( user_rst_n ),
    .received_func_lvl_rst_n                   ( cfg_received_func_lvl_rst_n ),
    .sys_rst_n                                 (~phy_rdy_n),
    .pl_rst_n                                  ( 1'b1 ),
    .dl_rst_n                                  ( 1'b1 ),
    .tl_rst_n                                  ( 1'b1 ),
    .cm_sticky_rst_n                           ( 1'b1 ),

    .func_lvl_rst_n                            ( func_lvl_rst_n ),
    .cm_rst_n                                  ( cm_rst_n ),
    .trn_rbar_hit                              ( trn_rbar_hit ),
    .trn_rd                                    ( trn_rd ),
    .trn_recrc_err                             ( trn_recrc_err ),
    .trn_reof                                  ( trn_reof ),
    .trn_rerrfwd                               ( trn_rerrfwd ),
    .trn_rrem                                  ( trn_rrem ),
    .trn_rsof                                  ( trn_rsof ),
    .trn_rsrc_dsc                              ( trn_rsrc_dsc ),
    .trn_rsrc_rdy                              ( trn_rsrc_rdy ),
    .trn_rdst_rdy                              ( trn_rdst_rdy ),
    .trn_rnp_ok                                ( rx_np_ok ),
    .trn_rnp_req                               ( rx_np_req ),
    .trn_rfcp_ret                              ( 1'b1 ),
    .trn_tbuf_av                               ( tx_buf_av ),
    .trn_tcfg_req                              ( tx_cfg_req ),
    .trn_tdllp_dst_rdy                         ( ),
    .trn_tdst_rdy                              ( trn_tdst_rdy ),
    .trn_terr_drop                             ( tx_err_drop ),
    .trn_tcfg_gnt                              ( trn_tcfg_gnt ),
    .trn_td                                    ( trn_td ),
    .trn_tdllp_data                            ( 32'b0 ),
    .trn_tdllp_src_rdy                         ( 1'b0 ),
    .trn_tecrc_gen                             ( trn_tecrc_gen ),
    .trn_teof                                  ( trn_teof ),
    .trn_terrfwd                               ( trn_terrfwd ),
    .trn_trem                                  ( trn_trem),
    .trn_tsof                                  ( trn_tsof ),
    .trn_tsrc_dsc                              ( trn_tsrc_dsc ),
    .trn_tsrc_rdy                              ( trn_tsrc_rdy ),
    .trn_tstr                                  ( trn_tstr ),

    .trn_fc_cpld                               ( fc_cpld ),
    .trn_fc_cplh                               ( fc_cplh ),
    .trn_fc_npd                                ( fc_npd ),
    .trn_fc_nph                                ( fc_nph ),
    .trn_fc_pd                                 ( fc_pd ),
    .trn_fc_ph                                 ( fc_ph ),
    .trn_fc_sel                                ( fc_sel ),

    .cfg_dev_id                                (cfg_dev_id),
    .cfg_vend_id                               (cfg_vend_id),
    .cfg_rev_id                                (cfg_rev_id),
    .cfg_subsys_id                             (cfg_subsys_id),
    .cfg_subsys_vend_id                        (cfg_subsys_vend_id),
    .cfg_pciecap_interrupt_msgnum              (cfg_pciecap_interrupt_msgnum),

    .cfg_bridge_serr_en                        (cfg_bridge_serr_en),

    .cfg_command_bus_master_enable             ( cfg_command_bus_master_enable ),
    .cfg_command_interrupt_disable             ( cfg_command_interrupt_disable ),
    .cfg_command_io_enable                     ( cfg_command_io_enable ),
    .cfg_command_mem_enable                    ( cfg_command_mem_enable ),
    .cfg_command_serr_en                       ( cfg_command_serr_en ),
    .cfg_dev_control_aux_power_en              ( cfg_dev_control_aux_power_en ),
    .cfg_dev_control_corr_err_reporting_en     ( cfg_dev_control_corr_err_reporting_en ),
    .cfg_dev_control_enable_ro                 ( cfg_dev_control_enable_ro ),
    .cfg_dev_control_ext_tag_en                ( cfg_dev_control_ext_tag_en ),
    .cfg_dev_control_fatal_err_reporting_en    ( cfg_dev_control_fatal_err_reporting_en ),
    .cfg_dev_control_max_payload               ( cfg_dev_control_max_payload ),
    .cfg_dev_control_max_read_req              ( cfg_dev_control_max_read_req ),
    .cfg_dev_control_non_fatal_reporting_en    ( cfg_dev_control_non_fatal_reporting_en ),
    .cfg_dev_control_no_snoop_en               ( cfg_dev_control_no_snoop_en ),
    .cfg_dev_control_phantom_en                ( cfg_dev_control_phantom_en ),
    .cfg_dev_control_ur_err_reporting_en       ( cfg_dev_control_ur_err_reporting_en ),
    .cfg_dev_control2_cpl_timeout_dis          ( cfg_dev_control2_cpl_timeout_dis ),
    .cfg_dev_control2_cpl_timeout_val          ( cfg_dev_control2_cpl_timeout_val ),
    .cfg_dev_control2_ari_forward_en           ( cfg_dev_control2_ari_forward_en),
    .cfg_dev_control2_atomic_requester_en      ( cfg_dev_control2_atomic_requester_en),
    .cfg_dev_control2_atomic_egress_block      ( cfg_dev_control2_atomic_egress_block),
    .cfg_dev_control2_ido_req_en               ( cfg_dev_control2_ido_req_en),
    .cfg_dev_control2_ido_cpl_en               ( cfg_dev_control2_ido_cpl_en),
    .cfg_dev_control2_ltr_en                   ( cfg_dev_control2_ltr_en),
    .cfg_dev_control2_tlp_prefix_block         ( cfg_dev_control2_tlp_prefix_block),
    .cfg_dev_status_corr_err_detected          ( cfg_dev_status_corr_err_detected ),
    .cfg_dev_status_fatal_err_detected         ( cfg_dev_status_fatal_err_detected ),
    .cfg_dev_status_non_fatal_err_detected     ( cfg_dev_status_non_fatal_err_detected ),
    .cfg_dev_status_ur_detected                ( cfg_dev_status_ur_detected ),

    .cfg_mgmt_do                               ( cfg_mgmt_do ),
    .cfg_err_aer_headerlog_set_n               ( cfg_err_aer_headerlog_set_n),
    .cfg_err_aer_headerlog                     ( cfg_err_aer_headerlog),
    .cfg_err_cpl_rdy_n                         ( cfg_err_cpl_rdy_n ),
    .cfg_interrupt_do                          ( cfg_interrupt_do ),
    .cfg_interrupt_mmenable                    ( cfg_interrupt_mmenable ),
    .cfg_interrupt_msienable                   ( cfg_interrupt_msienable ),
    .cfg_interrupt_msixenable                  ( cfg_interrupt_msixenable ),
    .cfg_interrupt_msixfm                      ( cfg_interrupt_msixfm ),
    .cfg_interrupt_rdy_n                       ( cfg_interrupt_rdy_n ),
    .cfg_link_control_rcb                      ( cfg_link_control_rcb ),
    .cfg_link_control_aspm_control             ( cfg_link_control_aspm_control ),
    .cfg_link_control_auto_bandwidth_int_en    ( cfg_link_control_auto_bandwidth_int_en ),
    .cfg_link_control_bandwidth_int_en         ( cfg_link_control_bandwidth_int_en ),
    .cfg_link_control_clock_pm_en              ( cfg_link_control_clock_pm_en ),
    .cfg_link_control_common_clock             ( cfg_link_control_common_clock ),
    .cfg_link_control_extended_sync            ( cfg_link_control_extended_sync ),
    .cfg_link_control_hw_auto_width_dis        ( cfg_link_control_hw_auto_width_dis ),
    .cfg_link_control_link_disable             ( cfg_link_control_link_disable ),
    .cfg_link_control_retrain_link             ( cfg_link_control_retrain_link ),
    .cfg_link_status_auto_bandwidth_status     ( cfg_link_status_auto_bandwidth_status ),
    .cfg_link_status_bandwidth_status          ( cfg_link_status_bandwidth_status ),
    .cfg_link_status_current_speed             ( cfg_link_status_current_speed ),
    .cfg_link_status_dll_active                ( cfg_link_status_dll_active ),
    .cfg_link_status_link_training             ( cfg_link_status_link_training ),
    .cfg_link_status_negotiated_width          ( cfg_link_status_negotiated_width),
    .cfg_msg_data                              ( cfg_msg_data ),
    .cfg_msg_received                          ( cfg_msg_received ),
    .cfg_msg_received_assert_int_a             ( cfg_msg_received_assert_int_a),
    .cfg_msg_received_assert_int_b             ( cfg_msg_received_assert_int_b),
    .cfg_msg_received_assert_int_c             ( cfg_msg_received_assert_int_c),
    .cfg_msg_received_assert_int_d             ( cfg_msg_received_assert_int_d),
    .cfg_msg_received_deassert_int_a           ( cfg_msg_received_deassert_int_a),
    .cfg_msg_received_deassert_int_b           ( cfg_msg_received_deassert_int_b),
    .cfg_msg_received_deassert_int_c           ( cfg_msg_received_deassert_int_c),
    .cfg_msg_received_deassert_int_d           ( cfg_msg_received_deassert_int_d),
    .cfg_msg_received_err_cor                  ( cfg_msg_received_err_cor),
    .cfg_msg_received_err_fatal                ( cfg_msg_received_err_fatal),
    .cfg_msg_received_err_non_fatal            ( cfg_msg_received_err_non_fatal),
    .cfg_msg_received_pm_as_nak                ( cfg_msg_received_pm_as_nak),
    .cfg_msg_received_pme_to                   ( cfg_msg_received_pme_to ),
    .cfg_msg_received_pme_to_ack               ( cfg_msg_received_pme_to_ack),
    .cfg_msg_received_pm_pme                   ( cfg_msg_received_pm_pme),
    .cfg_msg_received_setslotpowerlimit        ( cfg_msg_received_setslotpowerlimit),
    .cfg_msg_received_unlock                   ( cfg_msg_received_unlock),
    .cfg_pcie_link_state                       ( cfg_pcie_link_state ),
    .cfg_pmcsr_pme_en                          ( cfg_pmcsr_pme_en),
    .cfg_pmcsr_powerstate                      ( cfg_pmcsr_powerstate),
    .cfg_pmcsr_pme_status                      ( cfg_pmcsr_pme_status),
    .cfg_pm_rcv_as_req_l1_n                    ( cfg_pm_rcv_as_req_l1_n),
    .cfg_pm_rcv_enter_l1_n                     ( cfg_pm_rcv_enter_l1_n),
    .cfg_pm_rcv_enter_l23_n                    ( cfg_pm_rcv_enter_l23_n),

    .cfg_pm_rcv_req_ack_n                      ( cfg_pm_rcv_req_ack_n),
    .cfg_mgmt_rd_wr_done_n                     ( cfg_mgmt_rd_wr_done_n ),
    .cfg_slot_control_electromech_il_ctl_pulse (cfg_slot_control_electromech_il_ctl_pulse),
    .cfg_root_control_syserr_corr_err_en       ( cfg_root_control_syserr_corr_err_en),
    .cfg_root_control_syserr_non_fatal_err_en  ( cfg_root_control_syserr_non_fatal_err_en),
    .cfg_root_control_syserr_fatal_err_en      ( cfg_root_control_syserr_fatal_err_en),
    .cfg_root_control_pme_int_en               ( cfg_root_control_pme_int_en   ),
    .cfg_aer_ecrc_check_en                     ( cfg_aer_ecrc_check_en ),
    .cfg_aer_ecrc_gen_en                       ( cfg_aer_ecrc_gen_en ),
    .cfg_aer_rooterr_corr_err_reporting_en     ( cfg_aer_rooterr_corr_err_reporting_en),
    .cfg_aer_rooterr_non_fatal_err_reporting_en( cfg_aer_rooterr_non_fatal_err_reporting_en),
    .cfg_aer_rooterr_fatal_err_reporting_en    ( cfg_aer_rooterr_fatal_err_reporting_en),
    .cfg_aer_rooterr_corr_err_received         ( cfg_aer_rooterr_corr_err_received),
    .cfg_aer_rooterr_non_fatal_err_received    ( cfg_aer_rooterr_non_fatal_err_received),
    .cfg_aer_rooterr_fatal_err_received        ( cfg_aer_rooterr_fatal_err_received),
    .cfg_aer_interrupt_msgnum                  ( cfg_aer_interrupt_msgnum      ),
    .cfg_transaction                           ( cfg_transaction),
    .cfg_transaction_addr                      ( cfg_transaction_addr),
    .cfg_transaction_type                      ( cfg_transaction_type),
    .cfg_vc_tcvc_map                           ( cfg_vc_tcvc_map),
    .cfg_mgmt_byte_en_n                        ( cfg_mgmt_byte_en_n ),
    .cfg_mgmt_di                               ( cfg_mgmt_di ),
    .cfg_ds_bus_number                         ( cfg_ds_bus_number ),
    .cfg_ds_device_number                      ( cfg_ds_device_number ),
    .cfg_ds_function_number                    ( cfg_ds_function_number ),
    .cfg_dsn                                   ( cfg_dsn ),
    .cfg_mgmt_dwaddr                           ( cfg_mgmt_dwaddr ),
    .cfg_err_acs_n                             ( 1'b1 ),
    .cfg_err_cor_n                             ( cfg_err_cor_n ),
    .cfg_err_cpl_abort_n                       ( cfg_err_cpl_abort_n ),
    .cfg_err_cpl_timeout_n                     ( cfg_err_cpl_timeout_n ),
    .cfg_err_cpl_unexpect_n                    ( cfg_err_cpl_unexpect_n ),
    .cfg_err_ecrc_n                            ( cfg_err_ecrc_n ),
    .cfg_err_locked_n                          ( cfg_err_locked_n ),
    .cfg_err_posted_n                          ( cfg_err_posted_n ),
    .cfg_err_tlp_cpl_header                    ( cfg_err_tlp_cpl_header ),
    .cfg_err_ur_n                              ( cfg_err_ur_n ),
    .cfg_err_malformed_n                       ( cfg_err_malformed_n ),
    .cfg_err_poisoned_n                        ( cfg_err_poisoned_n),
    .cfg_err_atomic_egress_blocked_n           ( cfg_err_atomic_egress_blocked_n ),
    .cfg_err_mc_blocked_n                      ( cfg_err_mc_blocked_n  ),
    .cfg_err_internal_uncor_n                  ( cfg_err_internal_uncor_n      ),
    .cfg_err_internal_cor_n                    ( cfg_err_internal_cor_n ),
    .cfg_err_norecovery_n                      ( cfg_err_norecovery_n  ),

    .cfg_interrupt_assert_n                    ( cfg_interrupt_assert_n ),
    .cfg_interrupt_di                          ( cfg_interrupt_di ),
    .cfg_interrupt_n                           ( cfg_interrupt_n ),
    .cfg_interrupt_stat_n                      ( cfg_interrupt_stat_n),
    .cfg_pm_send_pme_to_n                      ( cfg_pm_send_pme_to_n ),
    .cfg_pm_turnoff_ok_n                       ( cfg_turnoff_ok_w ),
    .cfg_pm_wake_n                             ( cfg_pm_wake_n ),
    .cfg_pm_halt_aspm_l0s_n                    ( cfg_pm_halt_aspm_l0s_n ),
    .cfg_pm_halt_aspm_l1_n                     ( cfg_pm_halt_aspm_l1_n ),
    .cfg_pm_force_state_en_n                   ( cfg_pm_force_state_en_n ),
    .cfg_pm_force_state                        ( cfg_pm_force_state ),
    .cfg_force_mps                             ( cfg_force_mps ),
    .cfg_force_common_clock_off                ( cfg_force_common_clock_off ),
    .cfg_force_extended_sync_on                ( cfg_force_extended_sync_on ),
    .cfg_port_number                           ( cfg_port_number ),
    .cfg_mgmt_rd_en_n                          ( cfg_mgmt_rd_en_n ),
    .cfg_trn_pending_n                         ( ~cfg_trn_pending ),
    .cfg_mgmt_wr_en_n                          ( cfg_mgmt_wr_en_n ),
    .cfg_mgmt_wr_readonly_n                    ( cfg_mgmt_wr_readonly_n ),
    .cfg_mgmt_wr_rw1c_as_rw_n                  ( cfg_mgmt_wr_rw1c_as_rw_n ),

    .pl_initial_link_width                     ( pl_initial_link_width ),
    .pl_lane_reversal_mode                     ( pl_lane_reversal_mode ),
    .pl_link_gen2_cap                          ( pl_link_gen2_cap ),
    .pl_link_partner_gen2_supported            ( pl_link_partner_gen2_supported ),
    .pl_link_upcfg_cap                         ( pl_link_upcfg_cap ),
    .pl_ltssm_state                            ( pl_ltssm_state ),
    .pl_phy_lnk_up_n                           ( pl_phy_lnk_up_n ),
    .pl_received_hot_rst                       ( pl_received_hot_rst ),
    .pl_rx_pm_state                            ( pl_rx_pm_state ),
    .pl_sel_lnk_rate                           ( pl_sel_lnk_rate),
    .pl_sel_lnk_width                          ( pl_sel_lnk_width ),
    .pl_tx_pm_state                            ( pl_tx_pm_state ),
    .pl_directed_link_auton                    ( pl_directed_link_auton ),
    .pl_directed_link_change                   ( pl_directed_link_change ),
    .pl_directed_link_speed                    ( pl_directed_link_speed ),
    .pl_directed_link_width                    ( pl_directed_link_width ),
    .pl_downstream_deemph_source               ( pl_downstream_deemph_source ),
    .pl_upstream_prefer_deemph                 ( pl_upstream_prefer_deemph ),
    .pl_transmit_hot_rst                       ( pl_transmit_hot_rst ),
    .pl_directed_ltssm_new_vld                 ( pl_directed_ltssm_new_vld ),
    .pl_directed_ltssm_new                     ( pl_directed_ltssm_new ),
    .pl_directed_ltssm_stall                   ( pl_directed_ltssm_stall ),
    .pl_directed_change_done                   ( pl_directed_change_done ),

    .dbg_sclr_a                                ( dbg_sclr_a ),
    .dbg_sclr_b                                ( dbg_sclr_b ),
    .dbg_sclr_c                                ( dbg_sclr_c ),
    .dbg_sclr_d                                ( dbg_sclr_d ),
    .dbg_sclr_e                                ( dbg_sclr_e ),
    .dbg_sclr_f                                ( dbg_sclr_f ),
    .dbg_sclr_g                                ( dbg_sclr_g ),
    .dbg_sclr_h                                ( dbg_sclr_h ),
    .dbg_sclr_i                                ( dbg_sclr_i ),
    .dbg_sclr_j                                ( dbg_sclr_j ),
    .dbg_sclr_k                                ( dbg_sclr_k ),

    .dbg_vec_a                                 ( dbg_vec_a ),
    .dbg_vec_b                                 ( dbg_vec_b ),
    .dbg_vec_c                                 ( dbg_vec_c ),
    .pl_dbg_vec                                ( pl_dbg_vec ),
    .dbg_mode                                  ( dbg_mode ),
    .dbg_sub_mode                              ( dbg_sub_mode ),
    .pl_dbg_mode                               ( pl_dbg_mode ),

    .drp_do                                    ( drp_do ),
    .drp_rdy                                   ( drp_rdy ),
    .drp_clk                                   ( drp_clk ),
    .drp_addr                                  ( drp_addr ),
    .drp_en                                    ( drp_en ),
    .drp_di                                    ( drp_di ),
    .drp_we                                    ( drp_we ),

    .ll2_tlp_rcv                               ( 1'b0 ),
    .ll2_send_enter_l1                         ( 1'b0 ),
    .ll2_send_enter_l23                        ( 1'b0 ),
    .ll2_send_as_req_l1                        ( 1'b0 ),
    .ll2_send_pm_ack                           ( 1'b0 ),
    .ll2_suspend_now                           ( 1'b0 ),
    .ll2_tfc_init1_seq                         ( ),
    .ll2_tfc_init2_seq                         ( ),
    .ll2_suspend_ok                            ( ),
    .ll2_tx_idle                               ( ),
    .ll2_link_status                           ( ),
    .ll2_receiver_err                          ( ),
    .ll2_protocol_err                          ( ),
    .ll2_bad_tlp_err                           ( ),
    .ll2_bad_dllp_err                          ( ),
    .ll2_replay_ro_err                         ( ),
    .ll2_replay_to_err                         ( ),
    .tl2_ppm_suspend_req                       ( 1'b0 ),
    .tl2_aspm_suspend_credit_check             ( 1'b0 ),
    .tl2_ppm_suspend_ok                        ( ),
    .tl2_aspm_suspend_req                      ( ),
    .tl2_aspm_suspend_credit_check_ok          ( ),
    .tl2_err_hdr                               ( ),
    .tl2_err_malformed                         ( ),
    .tl2_err_rxoverflow                        ( ),
    .tl2_err_fcpe                              ( ),
    .pl2_directed_lstate                       ( 5'b0 ),
    .pl2_suspend_ok                            ( ),
    .pl2_recovery                              ( ),
    .pl2_rx_elec_idle                          ( ),
    .pl2_rx_pm_state                           ( ),
    .pl2_l0_req                                ( ),
    .pl2_link_up                               ( ),
    .pl2_receiver_err                          ( ),

    .trn_rdllp_data                            (trn_rdllp_data ),
    .trn_rdllp_src_rdy                         (trn_rdllp_src_rdy ),

    .pipe_clk                                  ( pipe_clk ),
    .user_clk2                                 ( user_clk2 ),
    .user_clk                                  ( user_clk ),
    .user_clk_prebuf                           ( 1'b0 ),
    .user_clk_prebuf_en                        ( 1'b0 ),

    .pipe_rx0_polarity                         ( pipe_rx0_polarity ),
    .pipe_rx1_polarity                         ( pipe_rx1_polarity ),
    .pipe_rx2_polarity                         ( pipe_rx2_polarity ),
    .pipe_rx3_polarity                         ( pipe_rx3_polarity ),
    .pipe_rx4_polarity                         ( pipe_rx4_polarity ),
    .pipe_rx5_polarity                         ( pipe_rx5_polarity ),
    .pipe_rx6_polarity                         ( pipe_rx6_polarity ),
    .pipe_rx7_polarity                         ( pipe_rx7_polarity ),
    .pipe_tx0_compliance                       ( pipe_tx0_compliance ),
    .pipe_tx1_compliance                       ( pipe_tx1_compliance ),
    .pipe_tx2_compliance                       ( pipe_tx2_compliance ),
    .pipe_tx3_compliance                       ( pipe_tx3_compliance ),
    .pipe_tx4_compliance                       ( pipe_tx4_compliance ),
    .pipe_tx5_compliance                       ( pipe_tx5_compliance ),
    .pipe_tx6_compliance                       ( pipe_tx6_compliance ),
    .pipe_tx7_compliance                       ( pipe_tx7_compliance ),
    .pipe_tx0_char_is_k                        ( pipe_tx0_char_is_k ),
    .pipe_tx1_char_is_k                        ( pipe_tx1_char_is_k ),
    .pipe_tx2_char_is_k                        ( pipe_tx2_char_is_k ),
    .pipe_tx3_char_is_k                        ( pipe_tx3_char_is_k ),
    .pipe_tx4_char_is_k                        ( pipe_tx4_char_is_k ),
    .pipe_tx5_char_is_k                        ( pipe_tx5_char_is_k ),
    .pipe_tx6_char_is_k                        ( pipe_tx6_char_is_k ),
    .pipe_tx7_char_is_k                        ( pipe_tx7_char_is_k ),
    .pipe_tx0_data                             ( pipe_tx0_data ),
    .pipe_tx1_data                             ( pipe_tx1_data ),
    .pipe_tx2_data                             ( pipe_tx2_data ),
    .pipe_tx3_data                             ( pipe_tx3_data ),
    .pipe_tx4_data                             ( pipe_tx4_data ),
    .pipe_tx5_data                             ( pipe_tx5_data ),
    .pipe_tx6_data                             ( pipe_tx6_data ),
    .pipe_tx7_data                             ( pipe_tx7_data ),
    .pipe_tx0_elec_idle                        ( pipe_tx0_elec_idle ),
    .pipe_tx1_elec_idle                        ( pipe_tx1_elec_idle ),
    .pipe_tx2_elec_idle                        ( pipe_tx2_elec_idle ),
    .pipe_tx3_elec_idle                        ( pipe_tx3_elec_idle ),
    .pipe_tx4_elec_idle                        ( pipe_tx4_elec_idle ),
    .pipe_tx5_elec_idle                        ( pipe_tx5_elec_idle ),
    .pipe_tx6_elec_idle                        ( pipe_tx6_elec_idle ),
    .pipe_tx7_elec_idle                        ( pipe_tx7_elec_idle ),
    .pipe_tx0_powerdown                        ( pipe_tx0_powerdown ),
    .pipe_tx1_powerdown                        ( pipe_tx1_powerdown ),
    .pipe_tx2_powerdown                        ( pipe_tx2_powerdown ),
    .pipe_tx3_powerdown                        ( pipe_tx3_powerdown ),
    .pipe_tx4_powerdown                        ( pipe_tx4_powerdown ),
    .pipe_tx5_powerdown                        ( pipe_tx5_powerdown ),
    .pipe_tx6_powerdown                        ( pipe_tx6_powerdown ),
    .pipe_tx7_powerdown                        ( pipe_tx7_powerdown ),

    .pipe_rx0_char_is_k                        ( pipe_rx0_char_is_k ),
    .pipe_rx1_char_is_k                        ( pipe_rx1_char_is_k ),
    .pipe_rx2_char_is_k                        ( pipe_rx2_char_is_k ),
    .pipe_rx3_char_is_k                        ( pipe_rx3_char_is_k ),
    .pipe_rx4_char_is_k                        ( pipe_rx4_char_is_k ),
    .pipe_rx5_char_is_k                        ( pipe_rx5_char_is_k ),
    .pipe_rx6_char_is_k                        ( pipe_rx6_char_is_k ),
    .pipe_rx7_char_is_k                        ( pipe_rx7_char_is_k ),
    .pipe_rx0_valid                            ( pipe_rx0_valid ),
    .pipe_rx1_valid                            ( pipe_rx1_valid ),
    .pipe_rx2_valid                            ( pipe_rx2_valid ),
    .pipe_rx3_valid                            ( pipe_rx3_valid ),
    .pipe_rx4_valid                            ( pipe_rx4_valid ),
    .pipe_rx5_valid                            ( pipe_rx5_valid ),
    .pipe_rx6_valid                            ( pipe_rx6_valid ),
    .pipe_rx7_valid                            ( pipe_rx7_valid ),
    .pipe_rx0_data                             ( pipe_rx0_data ),
    .pipe_rx1_data                             ( pipe_rx1_data ),
    .pipe_rx2_data                             ( pipe_rx2_data ),
    .pipe_rx3_data                             ( pipe_rx3_data ),
    .pipe_rx4_data                             ( pipe_rx4_data ),
    .pipe_rx5_data                             ( pipe_rx5_data ),
    .pipe_rx6_data                             ( pipe_rx6_data ),
    .pipe_rx7_data                             ( pipe_rx7_data ),
    .pipe_rx0_chanisaligned                    ( pipe_rx0_chanisaligned ),
    .pipe_rx1_chanisaligned                    ( pipe_rx1_chanisaligned ),
    .pipe_rx2_chanisaligned                    ( pipe_rx2_chanisaligned ),
    .pipe_rx3_chanisaligned                    ( pipe_rx3_chanisaligned ),
    .pipe_rx4_chanisaligned                    ( pipe_rx4_chanisaligned ),
    .pipe_rx5_chanisaligned                    ( pipe_rx5_chanisaligned ),
    .pipe_rx6_chanisaligned                    ( pipe_rx6_chanisaligned ),
    .pipe_rx7_chanisaligned                    ( pipe_rx7_chanisaligned ),
    .pipe_rx0_status                           ( pipe_rx0_status ),
    .pipe_rx1_status                           ( pipe_rx1_status ),
    .pipe_rx2_status                           ( pipe_rx2_status ),
    .pipe_rx3_status                           ( pipe_rx3_status ),
    .pipe_rx4_status                           ( pipe_rx4_status ),
    .pipe_rx5_status                           ( pipe_rx5_status ),
    .pipe_rx6_status                           ( pipe_rx6_status ),
    .pipe_rx7_status                           ( pipe_rx7_status ),
    .pipe_rx0_phy_status                       ( pipe_rx0_phy_status ),
    .pipe_rx1_phy_status                       ( pipe_rx1_phy_status ),
    .pipe_rx2_phy_status                       ( pipe_rx2_phy_status ),
    .pipe_rx3_phy_status                       ( pipe_rx3_phy_status ),
    .pipe_rx4_phy_status                       ( pipe_rx4_phy_status ),
    .pipe_rx5_phy_status                       ( pipe_rx5_phy_status ),
    .pipe_rx6_phy_status                       ( pipe_rx6_phy_status ),
    .pipe_rx7_phy_status                       ( pipe_rx7_phy_status ),
    .pipe_tx_deemph                            ( pipe_tx_deemph ),
    .pipe_tx_margin                            ( pipe_tx_margin ),
    .pipe_tx_reset                             ( pipe_tx_reset ),
    .pipe_tx_rcvr_det                          ( pipe_tx_rcvr_det ),
    .pipe_tx_rate                              ( pipe_tx_rate ),

    .pipe_rx0_elec_idle                        ( pipe_rx0_elec_idle ),
    .pipe_rx1_elec_idle                        ( pipe_rx1_elec_idle ),
    .pipe_rx2_elec_idle                        ( pipe_rx2_elec_idle ),
    .pipe_rx3_elec_idle                        ( pipe_rx3_elec_idle ),
    .pipe_rx4_elec_idle                        ( pipe_rx4_elec_idle ),
    .pipe_rx5_elec_idle                        ( pipe_rx5_elec_idle ),
    .pipe_rx6_elec_idle                        ( pipe_rx6_elec_idle ),
    .pipe_rx7_elec_idle                        ( pipe_rx7_elec_idle )
  );

  //------------------------------------------------------------------------------------------------------------------//
  // PIPE Interface PIPELINE Module                                                                                   //
  //------------------------------------------------------------------------------------------------------------------//
model_ap2_tst_pcie_pipe_pipeline # (

    .LINK_CAP_MAX_LINK_WIDTH ( LINK_CAP_MAX_LINK_WIDTH ),
    .PIPE_PIPELINE_STAGES    ( PIPE_PIPELINE_STAGES )

  )
  model_ap2_tst_pcie_pipe_pipeline_i (

    // Pipe Per-Link Signals
    .pipe_tx_rcvr_det_i       (pipe_tx_rcvr_det),
    .pipe_tx_reset_i          (1'b0), //MV?
    .pipe_tx_rate_i           (pipe_tx_rate),
    .pipe_tx_deemph_i         (pipe_tx_deemph),
    .pipe_tx_margin_i         (pipe_tx_margin),
    .pipe_tx_swing_i          (1'b0),

    .pipe_tx_rcvr_det_o       (pipe_tx_rcvr_det_gt),
    .pipe_tx_reset_o          ( ),
    .pipe_tx_rate_o           (pipe_tx_rate_gt),
    .pipe_tx_deemph_o         (pipe_tx_deemph_gt),
    .pipe_tx_margin_o         (pipe_tx_margin_gt),
    .pipe_tx_swing_o          ( ),

    // Pipe Per-Lane Signals - Lane 0

    .pipe_rx0_char_is_k_o     (pipe_rx0_char_is_k     ),
    .pipe_rx0_data_o          (pipe_rx0_data          ),
    .pipe_rx0_valid_o         (pipe_rx0_valid         ),
    .pipe_rx0_chanisaligned_o (pipe_rx0_chanisaligned ),
    .pipe_rx0_status_o        (pipe_rx0_status        ),
    .pipe_rx0_phy_status_o    (pipe_rx0_phy_status    ),
    .pipe_rx0_elec_idle_i     (pipe_rx0_elec_idle_gt  ),
    .pipe_rx0_polarity_i      (pipe_rx0_polarity      ),
    .pipe_tx0_compliance_i    (pipe_tx0_compliance    ),
    .pipe_tx0_char_is_k_i     (pipe_tx0_char_is_k     ),
    .pipe_tx0_data_i          (pipe_tx0_data          ),
    .pipe_tx0_elec_idle_i     (pipe_tx0_elec_idle     ),
    .pipe_tx0_powerdown_i     (pipe_tx0_powerdown     ),

    .pipe_rx0_char_is_k_i     (pipe_rx0_char_is_k_gt  ),
    .pipe_rx0_data_i          (pipe_rx0_data_gt       ),
    .pipe_rx0_valid_i         (pipe_rx0_valid_gt      ),
    .pipe_rx0_chanisaligned_i (pipe_rx0_chanisaligned_gt),
    .pipe_rx0_status_i        (pipe_rx0_status_gt     ),
    .pipe_rx0_phy_status_i    (pipe_rx0_phy_status_gt ),
    .pipe_rx0_elec_idle_o     (pipe_rx0_elec_idle     ),
    .pipe_rx0_polarity_o      (pipe_rx0_polarity_gt   ),
    .pipe_tx0_compliance_o    (pipe_tx0_compliance_gt ),
    .pipe_tx0_char_is_k_o     (pipe_tx0_char_is_k_gt  ),
    .pipe_tx0_data_o          (pipe_tx0_data_gt       ),
    .pipe_tx0_elec_idle_o     (pipe_tx0_elec_idle_gt  ),
    .pipe_tx0_powerdown_o     (pipe_tx0_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 1

    .pipe_rx1_char_is_k_o     (pipe_rx1_char_is_k     ),
    .pipe_rx1_data_o          (pipe_rx1_data          ),
    .pipe_rx1_valid_o         (pipe_rx1_valid         ),
    .pipe_rx1_chanisaligned_o (pipe_rx1_chanisaligned ),
    .pipe_rx1_status_o        (pipe_rx1_status        ),
    .pipe_rx1_phy_status_o    (pipe_rx1_phy_status    ),
    .pipe_rx1_elec_idle_i     (pipe_rx1_elec_idle_gt  ),
    .pipe_rx1_polarity_i      (pipe_rx1_polarity      ),
    .pipe_tx1_compliance_i    (pipe_tx1_compliance    ),
    .pipe_tx1_char_is_k_i     (pipe_tx1_char_is_k     ),
    .pipe_tx1_data_i          (pipe_tx1_data          ),
    .pipe_tx1_elec_idle_i     (pipe_tx1_elec_idle     ),
    .pipe_tx1_powerdown_i     (pipe_tx1_powerdown     ),

    .pipe_rx1_char_is_k_i     (pipe_rx1_char_is_k_gt  ),
    .pipe_rx1_data_i          (pipe_rx1_data_gt       ),
    .pipe_rx1_valid_i         (pipe_rx1_valid_gt      ),
    .pipe_rx1_chanisaligned_i (pipe_rx1_chanisaligned_gt),
    .pipe_rx1_status_i        (pipe_rx1_status_gt     ),
    .pipe_rx1_phy_status_i    (pipe_rx1_phy_status_gt ),
    .pipe_rx1_elec_idle_o     (pipe_rx1_elec_idle     ),
    .pipe_rx1_polarity_o      (pipe_rx1_polarity_gt   ),
    .pipe_tx1_compliance_o    (pipe_tx1_compliance_gt ),
    .pipe_tx1_char_is_k_o     (pipe_tx1_char_is_k_gt  ),
    .pipe_tx1_data_o          (pipe_tx1_data_gt       ),
    .pipe_tx1_elec_idle_o     (pipe_tx1_elec_idle_gt  ),
    .pipe_tx1_powerdown_o     (pipe_tx1_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 2

    .pipe_rx2_char_is_k_o     (pipe_rx2_char_is_k     ),
    .pipe_rx2_data_o          (pipe_rx2_data          ),
    .pipe_rx2_valid_o         (pipe_rx2_valid         ),
    .pipe_rx2_chanisaligned_o (pipe_rx2_chanisaligned ),
    .pipe_rx2_status_o        (pipe_rx2_status        ),
    .pipe_rx2_phy_status_o    (pipe_rx2_phy_status    ),
    .pipe_rx2_elec_idle_i     (pipe_rx2_elec_idle_gt  ),
    .pipe_rx2_polarity_i      (pipe_rx2_polarity      ),
    .pipe_tx2_compliance_i    (pipe_tx2_compliance    ),
    .pipe_tx2_char_is_k_i     (pipe_tx2_char_is_k     ),
    .pipe_tx2_data_i          (pipe_tx2_data          ),
    .pipe_tx2_elec_idle_i     (pipe_tx2_elec_idle     ),
    .pipe_tx2_powerdown_i     (pipe_tx2_powerdown     ),

    .pipe_rx2_char_is_k_i     (pipe_rx2_char_is_k_gt  ),
    .pipe_rx2_data_i          (pipe_rx2_data_gt       ),
    .pipe_rx2_valid_i         (pipe_rx2_valid_gt      ),
    .pipe_rx2_chanisaligned_i (pipe_rx2_chanisaligned_gt),
    .pipe_rx2_status_i        (pipe_rx2_status_gt     ),
    .pipe_rx2_phy_status_i    (pipe_rx2_phy_status_gt ),
    .pipe_rx2_elec_idle_o     (pipe_rx2_elec_idle     ),
    .pipe_rx2_polarity_o      (pipe_rx2_polarity_gt   ),
    .pipe_tx2_compliance_o    (pipe_tx2_compliance_gt ),
    .pipe_tx2_char_is_k_o     (pipe_tx2_char_is_k_gt  ),
    .pipe_tx2_data_o          (pipe_tx2_data_gt       ),
    .pipe_tx2_elec_idle_o     (pipe_tx2_elec_idle_gt  ),
    .pipe_tx2_powerdown_o     (pipe_tx2_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 3

    .pipe_rx3_char_is_k_o     (pipe_rx3_char_is_k     ),
    .pipe_rx3_data_o          (pipe_rx3_data          ),
    .pipe_rx3_valid_o         (pipe_rx3_valid         ),
    .pipe_rx3_chanisaligned_o (pipe_rx3_chanisaligned ),
    .pipe_rx3_status_o        (pipe_rx3_status        ),
    .pipe_rx3_phy_status_o    (pipe_rx3_phy_status    ),
    .pipe_rx3_elec_idle_i     (pipe_rx3_elec_idle_gt  ),
    .pipe_rx3_polarity_i      (pipe_rx3_polarity      ),
    .pipe_tx3_compliance_i    (pipe_tx3_compliance    ),
    .pipe_tx3_char_is_k_i     (pipe_tx3_char_is_k     ),
    .pipe_tx3_data_i          (pipe_tx3_data          ),
    .pipe_tx3_elec_idle_i     (pipe_tx3_elec_idle     ),
    .pipe_tx3_powerdown_i     (pipe_tx3_powerdown     ),

    .pipe_rx3_char_is_k_i     (pipe_rx3_char_is_k_gt  ),
    .pipe_rx3_data_i          (pipe_rx3_data_gt       ),
    .pipe_rx3_valid_i         (pipe_rx3_valid_gt      ),
    .pipe_rx3_chanisaligned_i (pipe_rx3_chanisaligned_gt),
    .pipe_rx3_status_i        (pipe_rx3_status_gt     ),
    .pipe_rx3_phy_status_i    (pipe_rx3_phy_status_gt ),
    .pipe_rx3_elec_idle_o     (pipe_rx3_elec_idle     ),
    .pipe_rx3_polarity_o      (pipe_rx3_polarity_gt   ),
    .pipe_tx3_compliance_o    (pipe_tx3_compliance_gt ),
    .pipe_tx3_char_is_k_o     (pipe_tx3_char_is_k_gt  ),
    .pipe_tx3_data_o          (pipe_tx3_data_gt       ),
    .pipe_tx3_elec_idle_o     (pipe_tx3_elec_idle_gt  ),
    .pipe_tx3_powerdown_o     (pipe_tx3_powerdown_gt  ),

     // Pipe Per-Lane Signals - Lane 4

    .pipe_rx4_char_is_k_o     (pipe_rx4_char_is_k     ),
    .pipe_rx4_data_o          (pipe_rx4_data          ),
    .pipe_rx4_valid_o         (pipe_rx4_valid         ),
    .pipe_rx4_chanisaligned_o (pipe_rx4_chanisaligned ),
    .pipe_rx4_status_o        (pipe_rx4_status        ),
    .pipe_rx4_phy_status_o    (pipe_rx4_phy_status    ),
    .pipe_rx4_elec_idle_i     (pipe_rx4_elec_idle_gt  ),
    .pipe_rx4_polarity_i      (pipe_rx4_polarity      ),
    .pipe_tx4_compliance_i    (pipe_tx4_compliance    ),
    .pipe_tx4_char_is_k_i     (pipe_tx4_char_is_k     ),
    .pipe_tx4_data_i          (pipe_tx4_data          ),
    .pipe_tx4_elec_idle_i     (pipe_tx4_elec_idle     ),
    .pipe_tx4_powerdown_i     (pipe_tx4_powerdown     ),
    .pipe_rx4_char_is_k_i     (pipe_rx4_char_is_k_gt  ),
    .pipe_rx4_data_i          (pipe_rx4_data_gt       ),
    .pipe_rx4_valid_i         (pipe_rx4_valid_gt      ),
    .pipe_rx4_chanisaligned_i (pipe_rx4_chanisaligned_gt),
    .pipe_rx4_status_i        (pipe_rx4_status_gt     ),
    .pipe_rx4_phy_status_i    (pipe_rx4_phy_status_gt ),
    .pipe_rx4_elec_idle_o     (pipe_rx4_elec_idle     ),
    .pipe_rx4_polarity_o      (pipe_rx4_polarity_gt   ),
    .pipe_tx4_compliance_o    (pipe_tx4_compliance_gt ),
    .pipe_tx4_char_is_k_o     (pipe_tx4_char_is_k_gt  ),
    .pipe_tx4_data_o          (pipe_tx4_data_gt       ),
    .pipe_tx4_elec_idle_o     (pipe_tx4_elec_idle_gt  ),
    .pipe_tx4_powerdown_o     (pipe_tx4_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 5

    .pipe_rx5_char_is_k_o     (pipe_rx5_char_is_k     ),
    .pipe_rx5_data_o          (pipe_rx5_data          ),
    .pipe_rx5_valid_o         (pipe_rx5_valid         ),
    .pipe_rx5_chanisaligned_o (pipe_rx5_chanisaligned ),
    .pipe_rx5_status_o        (pipe_rx5_status        ),
    .pipe_rx5_phy_status_o    (pipe_rx5_phy_status    ),
    .pipe_rx5_elec_idle_i     (pipe_rx5_elec_idle_gt  ),
    .pipe_rx5_polarity_i      (pipe_rx5_polarity      ),
    .pipe_tx5_compliance_i    (pipe_tx5_compliance    ),
    .pipe_tx5_char_is_k_i     (pipe_tx5_char_is_k     ),
    .pipe_tx5_data_i          (pipe_tx5_data          ),
    .pipe_tx5_elec_idle_i     (pipe_tx5_elec_idle     ),
    .pipe_tx5_powerdown_i     (pipe_tx5_powerdown     ),
    .pipe_rx5_char_is_k_i     (pipe_rx5_char_is_k_gt  ),
    .pipe_rx5_data_i          (pipe_rx5_data_gt       ),
    .pipe_rx5_valid_i         (pipe_rx5_valid_gt      ),
    .pipe_rx5_chanisaligned_i (pipe_rx5_chanisaligned_gt),
    .pipe_rx5_status_i        (pipe_rx5_status_gt     ),
    .pipe_rx5_phy_status_i    (pipe_rx5_phy_status_gt ),
    .pipe_rx5_elec_idle_o     (pipe_rx5_elec_idle     ),
    .pipe_rx5_polarity_o      (pipe_rx5_polarity_gt   ),
    .pipe_tx5_compliance_o    (pipe_tx5_compliance_gt ),
    .pipe_tx5_char_is_k_o     (pipe_tx5_char_is_k_gt  ),
    .pipe_tx5_data_o          (pipe_tx5_data_gt       ),
    .pipe_tx5_elec_idle_o     (pipe_tx5_elec_idle_gt  ),
    .pipe_tx5_powerdown_o     (pipe_tx5_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 6

    .pipe_rx6_char_is_k_o     (pipe_rx6_char_is_k     ),
    .pipe_rx6_data_o          (pipe_rx6_data          ),
    .pipe_rx6_valid_o         (pipe_rx6_valid         ),
    .pipe_rx6_chanisaligned_o (pipe_rx6_chanisaligned ),
    .pipe_rx6_status_o        (pipe_rx6_status        ),
    .pipe_rx6_phy_status_o    (pipe_rx6_phy_status    ),
    .pipe_rx6_elec_idle_i     (pipe_rx6_elec_idle_gt  ),
    .pipe_rx6_polarity_i      (pipe_rx6_polarity      ),
    .pipe_tx6_compliance_i    (pipe_tx6_compliance    ),
    .pipe_tx6_char_is_k_i     (pipe_tx6_char_is_k     ),
    .pipe_tx6_data_i          (pipe_tx6_data          ),
    .pipe_tx6_elec_idle_i     (pipe_tx6_elec_idle     ),
    .pipe_tx6_powerdown_i     (pipe_tx6_powerdown     ),
    .pipe_rx6_char_is_k_i     (pipe_rx6_char_is_k_gt  ),
    .pipe_rx6_data_i          (pipe_rx6_data_gt       ),
    .pipe_rx6_valid_i         (pipe_rx6_valid_gt      ),
    .pipe_rx6_chanisaligned_i (pipe_rx6_chanisaligned_gt),
    .pipe_rx6_status_i        (pipe_rx6_status_gt     ),
    .pipe_rx6_phy_status_i    (pipe_rx6_phy_status_gt ),
    .pipe_rx6_elec_idle_o     (pipe_rx6_elec_idle     ),
    .pipe_rx6_polarity_o      (pipe_rx6_polarity_gt   ),
    .pipe_tx6_compliance_o    (pipe_tx6_compliance_gt ),
    .pipe_tx6_char_is_k_o     (pipe_tx6_char_is_k_gt  ),
    .pipe_tx6_data_o          (pipe_tx6_data_gt       ),
    .pipe_tx6_elec_idle_o     (pipe_tx6_elec_idle_gt  ),
    .pipe_tx6_powerdown_o     (pipe_tx6_powerdown_gt  ),

    // Pipe Per-Lane Signals - Lane 7

    .pipe_rx7_char_is_k_o     (pipe_rx7_char_is_k     ),
    .pipe_rx7_data_o          (pipe_rx7_data          ),
    .pipe_rx7_valid_o         (pipe_rx7_valid         ),
    .pipe_rx7_chanisaligned_o (pipe_rx7_chanisaligned ),
    .pipe_rx7_status_o        (pipe_rx7_status        ),
    .pipe_rx7_phy_status_o    (pipe_rx7_phy_status    ),
    .pipe_rx7_elec_idle_i     (pipe_rx7_elec_idle_gt  ),
    .pipe_rx7_polarity_i      (pipe_rx7_polarity      ),
    .pipe_tx7_compliance_i    (pipe_tx7_compliance    ),
    .pipe_tx7_char_is_k_i     (pipe_tx7_char_is_k     ),
    .pipe_tx7_data_i          (pipe_tx7_data          ),
    .pipe_tx7_elec_idle_i     (pipe_tx7_elec_idle     ),
    .pipe_tx7_powerdown_i     (pipe_tx7_powerdown     ),
    .pipe_rx7_char_is_k_i     (pipe_rx7_char_is_k_gt  ),
    .pipe_rx7_data_i          (pipe_rx7_data_gt       ),
    .pipe_rx7_valid_i         (pipe_rx7_valid_gt      ),
    .pipe_rx7_chanisaligned_i (pipe_rx7_chanisaligned_gt),
    .pipe_rx7_status_i        (pipe_rx7_status_gt     ),
    .pipe_rx7_phy_status_i    (pipe_rx7_phy_status_gt ),
    .pipe_rx7_elec_idle_o     (pipe_rx7_elec_idle     ),
    .pipe_rx7_polarity_o      (pipe_rx7_polarity_gt   ),
    .pipe_tx7_compliance_o    (pipe_tx7_compliance_gt ),
    .pipe_tx7_char_is_k_o     (pipe_tx7_char_is_k_gt  ),
    .pipe_tx7_data_o          (pipe_tx7_data_gt       ),
    .pipe_tx7_elec_idle_o     (pipe_tx7_elec_idle_gt  ),
    .pipe_tx7_powerdown_o     (pipe_tx7_powerdown_gt  ),

    // Non PIPE signals
    .pipe_clk                 (pipe_clk               ),
    .rst_n                    (phy_rdy_n              )
  );



endmodule




`timescale 1ns/1ps
module model_ap2_tst_axi_basic_top #(
  parameter C_DATA_WIDTH  = 128,          // RX/TX interface data width
  parameter C_FAMILY      = "X7",         // Targeted FPGA family
  parameter C_ROOT_PORT   = "FALSE",      // PCIe block is in root port mode
  parameter C_PM_PRIORITY = "FALSE",      // Disable TX packet boundary thrtl
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter REM_WIDTH  = (C_DATA_WIDTH == 128) ? 2 : 1, // trem/rrem width
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8               // KEEP width
  ) (
  //---------------------------------------------//
  // User Design I/O                             //
  //---------------------------------------------//

  // AXI TX
  //-----------
  input   [C_DATA_WIDTH-1:0] s_axis_tx_tdata,        // TX data from user
  input                      s_axis_tx_tvalid,       // TX data is valid
  output                     s_axis_tx_tready,       // TX ready for data
  input     [KEEP_WIDTH-1:0] s_axis_tx_tkeep,        // TX strobe byte enables
  input                      s_axis_tx_tlast,        // TX data is last
  input                [3:0] s_axis_tx_tuser,        // TX user signals

  // AXI RX
  //-----------
  output  [C_DATA_WIDTH-1:0] m_axis_rx_tdata,        // RX data to user
  output                     m_axis_rx_tvalid,       // RX data is valid
  input                      m_axis_rx_tready,       // RX ready for data
  output    [KEEP_WIDTH-1:0] m_axis_rx_tkeep,        // RX strobe byte enables
  output                     m_axis_rx_tlast,        // RX data is last
  output              [21:0] m_axis_rx_tuser,        // RX user signals

  // User Misc.
  //-----------
  input                      user_turnoff_ok,        // Turnoff OK from user
  input                      user_tcfg_gnt,          // Send cfg OK from user

  //---------------------------------------------//
  // PCIe Block I/O                              //
  //---------------------------------------------//

  // TRN TX
  //-----------
  output [C_DATA_WIDTH-1:0] trn_td,                  // TX data from block
  output                    trn_tsof,                // TX start of packet
  output                    trn_teof,                // TX end of packet
  output                    trn_tsrc_rdy,            // TX source ready
  input                     trn_tdst_rdy,            // TX destination ready
  output                    trn_tsrc_dsc,            // TX source discontinue
  output    [REM_WIDTH-1:0] trn_trem,                // TX remainder
  output                    trn_terrfwd,             // TX error forward
  output                    trn_tstr,                // TX streaming enable
  input               [5:0] trn_tbuf_av,             // TX buffers available
  output                    trn_tecrc_gen,           // TX ECRC generate

  // TRN RX
  //-----------
  input  [127:0] trn_rd,                  // RX data from block
  input                     trn_rsof,                // RX start of packet
  input                     trn_reof,                // RX end of packet
  input                     trn_rsrc_rdy,            // RX source ready
  output                    trn_rdst_rdy,            // RX destination ready
  input                     trn_rsrc_dsc,            // RX source discontinue
  input     [1:0] trn_rrem,                // RX remainder
  input                     trn_rerrfwd,             // RX error forward
  input               [6:0] trn_rbar_hit,            // RX BAR hit
  input                     trn_recrc_err,           // RX ECRC error

  // TRN Misc.
  //-----------
  input                     trn_tcfg_req,            // TX config request
  output                    trn_tcfg_gnt,            // RX config grant
  input                     trn_lnk_up,              // PCIe link up

  // 7 Series/Virtex6 PM
  //-----------
  input               [2:0] cfg_pcie_link_state,     // Encoded PCIe link state

  // Virtex6 PM
  //-----------
  input                     cfg_pm_send_pme_to,      // PM send PME turnoff msg
  input               [1:0] cfg_pmcsr_powerstate,    // PMCSR power state
  input              [31:0] trn_rdllp_data,          // RX DLLP data
  input                     trn_rdllp_src_rdy,       // RX DLLP source ready

  // Virtex6/Spartan6 PM
  //-----------
  input                     cfg_to_turnoff,          // Turnoff request
  output                    cfg_turnoff_ok,          // Turnoff grant

  // System
  //-----------
  output              [2:0] np_counter,              // Non-posted counter
  input                     user_clk,                // user clock from block
  input                     user_rst                 // user reset from block
);


//---------------------------------------------//
// RX Data Pipeline                            //
//---------------------------------------------//

model_ap2_tst_axi_basic_rx #(
  .C_DATA_WIDTH( C_DATA_WIDTH ),
  .C_FAMILY( C_FAMILY ),

  .TCQ( TCQ ),
  .REM_WIDTH( REM_WIDTH ),
  .KEEP_WIDTH( KEEP_WIDTH )
) model_ap2_tst_rx_inst (

  // Outgoing AXI TX
  //-----------
  .m_axis_rx_tdata( m_axis_rx_tdata ),
  .m_axis_rx_tvalid( m_axis_rx_tvalid ),
  .m_axis_rx_tready( m_axis_rx_tready ),
  .m_axis_rx_tkeep( m_axis_rx_tkeep ),
  .m_axis_rx_tlast( m_axis_rx_tlast ),
  .m_axis_rx_tuser( m_axis_rx_tuser ),

  // Incoming TRN RX
  //-----------
  .trn_rd( trn_rd[C_DATA_WIDTH-1:0] ),
  .trn_rsof( trn_rsof ),
  .trn_reof( trn_reof ),
  .trn_rsrc_rdy( trn_rsrc_rdy ),
  .trn_rdst_rdy( trn_rdst_rdy ),
  .trn_rsrc_dsc( trn_rsrc_dsc ),
  .trn_rrem( trn_rrem[REM_WIDTH-1:0] ),
  .trn_rerrfwd( trn_rerrfwd ),
  .trn_rbar_hit( trn_rbar_hit ),
  .trn_recrc_err( trn_recrc_err ),

  // System
  //-----------
  .np_counter( np_counter ),
  .user_clk( user_clk ),
  .user_rst( user_rst )
);



//---------------------------------------------//
// TX Data Pipeline                            //
//---------------------------------------------//

model_ap2_tst_axi_basic_tx #(
  .C_DATA_WIDTH( C_DATA_WIDTH ),
  .C_FAMILY( C_FAMILY ),
  .C_ROOT_PORT( C_ROOT_PORT ),
  .C_PM_PRIORITY( C_PM_PRIORITY ),

  .TCQ( TCQ ),
  .REM_WIDTH( REM_WIDTH ),
  .KEEP_WIDTH( KEEP_WIDTH )
) model_ap2_tst_tx_inst (

  // Incoming AXI RX
  //-----------
  .s_axis_tx_tdata( s_axis_tx_tdata ),
  .s_axis_tx_tvalid( s_axis_tx_tvalid ),
  .s_axis_tx_tready( s_axis_tx_tready ),
  .s_axis_tx_tkeep( s_axis_tx_tkeep ),
  .s_axis_tx_tlast( s_axis_tx_tlast ),
  .s_axis_tx_tuser( s_axis_tx_tuser ),

  // User Misc.
  //-----------
  .user_turnoff_ok( user_turnoff_ok ),
  .user_tcfg_gnt( user_tcfg_gnt ),

  // Outgoing TRN TX
  //-----------
  .trn_td( trn_td ),
  .trn_tsof( trn_tsof ),
  .trn_teof( trn_teof ),
  .trn_tsrc_rdy( trn_tsrc_rdy ),
  .trn_tdst_rdy( trn_tdst_rdy ),
  .trn_tsrc_dsc( trn_tsrc_dsc ),
  .trn_trem( trn_trem ),
  .trn_terrfwd( trn_terrfwd ),
  .trn_tstr( trn_tstr ),
  .trn_tbuf_av( trn_tbuf_av ),
  .trn_tecrc_gen( trn_tecrc_gen ),

  // TRN Misc.
  //-----------
  .trn_tcfg_req( trn_tcfg_req ),
  .trn_tcfg_gnt( trn_tcfg_gnt ),
  .trn_lnk_up( trn_lnk_up ),

  // 7 Series/Virtex6 PM
  //-----------
  .cfg_pcie_link_state( cfg_pcie_link_state ),

  // Virtex6 PM
  //-----------
  .cfg_pm_send_pme_to( cfg_pm_send_pme_to ),
  .cfg_pmcsr_powerstate( cfg_pmcsr_powerstate ),
  .trn_rdllp_data( trn_rdllp_data ),
  .trn_rdllp_src_rdy( trn_rdllp_src_rdy ),

  // Spartan6 PM
  //-----------
  .cfg_to_turnoff( cfg_to_turnoff ),
  .cfg_turnoff_ok( cfg_turnoff_ok ),

  // System
  //-----------
  .user_clk( user_clk ),
  .user_rst( user_rst )
);

endmodule


`timescale 1ns/1ps
module model_ap2_tst_axi_basic_rx #(
  parameter C_DATA_WIDTH  = 128,          // RX/TX interface data width
  parameter C_FAMILY      = "X7",         // Targeted FPGA family
  parameter C_ROOT_PORT   = "FALSE",      // PCIe block is in root port mode
  parameter C_PM_PRIORITY = "FALSE",      // Disable TX packet boundary thrtl
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter REM_WIDTH  = (C_DATA_WIDTH == 128) ? 2 : 1, // trem/rrem width
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8               // KEEP width
  ) (
  //---------------------------------------------//
  // User Design I/O                             //
  //---------------------------------------------//

  // AXI RX
  //-----------
  output  [C_DATA_WIDTH-1:0] m_axis_rx_tdata,        // RX data to user
  output                     m_axis_rx_tvalid,       // RX data is valid
  input                      m_axis_rx_tready,       // RX ready for data
  output    [KEEP_WIDTH-1:0] m_axis_rx_tkeep,        // RX strobe byte enables
  output                     m_axis_rx_tlast,        // RX data is last
  output              [21:0] m_axis_rx_tuser,        // RX user signals

  //---------------------------------------------//
  // PCIe Block I/O                              //
  //---------------------------------------------//

  // TRN RX
  //-----------
  input  [C_DATA_WIDTH-1:0] trn_rd,                  // RX data from block
  input                     trn_rsof,                // RX start of packet
  input                     trn_reof,                // RX end of packet
  input                     trn_rsrc_rdy,            // RX source ready
  output                    trn_rdst_rdy,            // RX destination ready
  input                     trn_rsrc_dsc,            // RX source discontinue
  input     [REM_WIDTH-1:0] trn_rrem,                // RX remainder
  input                     trn_rerrfwd,             // RX error forward
  input               [6:0] trn_rbar_hit,            // RX BAR hit
  input                     trn_recrc_err,           // RX ECRC error

  // System
  //-----------
  output              [2:0] np_counter,              // Non-posted counter
  input                     user_clk,                // user clock from block
  input                     user_rst                 // user reset from block
);


// Wires
wire                  null_rx_tvalid;
wire                  null_rx_tlast;
wire [KEEP_WIDTH-1:0] null_rx_tkeep;
wire                  null_rdst_rdy;
wire            [4:0] null_is_eof;

//---------------------------------------------//
// RX Data Pipeline                            //
//---------------------------------------------//

model_ap2_tst_axi_basic_rx_pipeline #(
  .C_DATA_WIDTH( C_DATA_WIDTH ),
  .C_FAMILY( C_FAMILY ),
  .TCQ( TCQ ),

  .REM_WIDTH( REM_WIDTH ),
  .KEEP_WIDTH( KEEP_WIDTH )

) model_ap2_tst_rx_pipeline_inst (

  // Outgoing AXI TX
  //-----------
  .m_axis_rx_tdata( m_axis_rx_tdata ),
  .m_axis_rx_tvalid( m_axis_rx_tvalid ),
  .m_axis_rx_tready( m_axis_rx_tready ),
  .m_axis_rx_tkeep( m_axis_rx_tkeep ),
  .m_axis_rx_tlast( m_axis_rx_tlast ),
  .m_axis_rx_tuser( m_axis_rx_tuser ),

  // Incoming TRN RX
  //-----------
  .trn_rd( trn_rd ),
  .trn_rsof( trn_rsof ),
  .trn_reof( trn_reof ),
  .trn_rsrc_rdy( trn_rsrc_rdy ),
  .trn_rdst_rdy( trn_rdst_rdy ),
  .trn_rsrc_dsc( trn_rsrc_dsc ),
  .trn_rrem( trn_rrem ),
  .trn_rerrfwd( trn_rerrfwd ),
  .trn_rbar_hit( trn_rbar_hit ),
  .trn_recrc_err( trn_recrc_err ),

  // Null Inputs
  //-----------
  .null_rx_tvalid( null_rx_tvalid ),
  .null_rx_tlast( null_rx_tlast ),
  .null_rx_tkeep( null_rx_tkeep ),
  .null_rdst_rdy( null_rdst_rdy ),
  .null_is_eof( null_is_eof ),

  // System
  //-----------
  .np_counter( np_counter ),
  .user_clk( user_clk ),
  .user_rst( user_rst )
);


 //---------------------------------------------//
 // RX Null Packet Generator                    //
 //---------------------------------------------//

model_ap2_tst_axi_basic_rx_null_gen #(
  .C_DATA_WIDTH( C_DATA_WIDTH ),
  .TCQ( TCQ ),

  .KEEP_WIDTH( KEEP_WIDTH )

 ) model_ap2_tst_rx_null_gen_inst (

  // Inputs
  //-----------
  .m_axis_rx_tdata( m_axis_rx_tdata ),
  .m_axis_rx_tvalid( m_axis_rx_tvalid ),
  .m_axis_rx_tready( m_axis_rx_tready ),
  .m_axis_rx_tlast( m_axis_rx_tlast ),
  .m_axis_rx_tuser( m_axis_rx_tuser ),

  // Null Outputs
  //-----------
  .null_rx_tvalid( null_rx_tvalid ),
  .null_rx_tlast( null_rx_tlast ),
  .null_rx_tkeep( null_rx_tkeep ),
  .null_rdst_rdy( null_rdst_rdy ),
  .null_is_eof( null_is_eof ),

  // System
  //-----------
  .user_clk( user_clk ),
  .user_rst( user_rst )
 );

endmodule



`timescale 1ns/1ps
module model_ap2_tst_axi_basic_rx_pipeline #(
  parameter C_DATA_WIDTH = 128,           // RX/TX interface data width
  parameter C_FAMILY     = "X7",          // Targeted FPGA family
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter REM_WIDTH  = (C_DATA_WIDTH == 128) ? 2 : 1, // trem/rrem width
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8               // KEEP width
  ) (

  // AXI RX
  //-----------
  output reg [C_DATA_WIDTH-1:0] m_axis_rx_tdata,     // RX data to user
  output reg                    m_axis_rx_tvalid,    // RX data is valid
  input                         m_axis_rx_tready,    // RX ready for data
  output       [KEEP_WIDTH-1:0] m_axis_rx_tkeep,     // RX strobe byte enables
  output                        m_axis_rx_tlast,     // RX data is last
  output reg             [21:0] m_axis_rx_tuser,     // RX user signals

  // TRN RX
  //-----------
  input      [C_DATA_WIDTH-1:0] trn_rd,              // RX data from block
  input                         trn_rsof,            // RX start of packet
  input                         trn_reof,            // RX end of packet
  input                         trn_rsrc_rdy,        // RX source ready
  output reg                    trn_rdst_rdy,        // RX destination ready
  input                         trn_rsrc_dsc,        // RX source discontinue
  input         [REM_WIDTH-1:0] trn_rrem,            // RX remainder
  input                         trn_rerrfwd,         // RX error forward
  input                   [6:0] trn_rbar_hit,        // RX BAR hit
  input                         trn_recrc_err,       // RX ECRC error

  // Null Inputs
  //-----------
  input                         null_rx_tvalid,      // NULL generated tvalid
  input                         null_rx_tlast,       // NULL generated tlast
  input        [KEEP_WIDTH-1:0] null_rx_tkeep,       // NULL generated tkeep
  input                         null_rdst_rdy,       // NULL generated rdst_rdy
  input                   [4:0] null_is_eof,         // NULL generated is_eof

  // System
  //-----------
  output                  [2:0] np_counter,          // Non-posted counter
  input                         user_clk,            // user clock from block
  input                         user_rst             // user reset from block
);


// Wires and regs for creating AXI signals
wire              [4:0] is_sof;
wire              [4:0] is_sof_prev;

wire              [4:0] is_eof;
wire              [4:0] is_eof_prev;

reg    [KEEP_WIDTH-1:0] reg_tkeep;
wire   [KEEP_WIDTH-1:0] tkeep;
wire   [KEEP_WIDTH-1:0] tkeep_prev;

reg                     reg_tlast;
wire                    rsrc_rdy_filtered;

// Wires and regs for previous value buffer
wire [C_DATA_WIDTH-1:0] trn_rd_DW_swapped;
reg  [C_DATA_WIDTH-1:0] trn_rd_prev;

wire                    data_hold;
reg                     data_prev;

reg                     trn_reof_prev;
reg     [REM_WIDTH-1:0] trn_rrem_prev;
reg                     trn_rsrc_rdy_prev;
reg                     trn_rsrc_dsc_prev;
reg                     trn_rsof_prev;
reg               [6:0] trn_rbar_hit_prev;
reg                     trn_rerrfwd_prev;
reg                     trn_recrc_err_prev;

// Null packet handling signals
reg                     null_mux_sel;
reg                     trn_in_packet;
wire                    dsc_flag;
wire                    dsc_detect;
reg                     reg_dsc_detect;
reg                     trn_rsrc_dsc_d;


// Create "filtered" version of rsrc_rdy, where discontinued SOFs are removed.
assign rsrc_rdy_filtered = trn_rsrc_rdy &&
                                 (trn_in_packet || (trn_rsof && !trn_rsrc_dsc));

//----------------------------------------------------------------------------//
// Previous value buffer                                                      //
// ---------------------                                                      //
// We are inserting a pipeline stage in between TRN and AXI, which causes     //
// some issues with handshaking signals m_axis_rx_tready/trn_rdst_rdy. The    //
// added cycle of latency in the path causes the user design to fall behind   //
// the TRN interface whenever it throttles.                                   //
//                                                                            //
// To avoid loss of data, we must keep the previous value of all trn_r*       //
// signals in case the user throttles.                                        //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    trn_rd_prev        <= #TCQ {C_DATA_WIDTH{1'b0}};
    trn_rsof_prev      <= #TCQ 1'b0;
    trn_rrem_prev      <= #TCQ {REM_WIDTH{1'b0}};
    trn_rsrc_rdy_prev  <= #TCQ 1'b0;
    trn_rbar_hit_prev  <= #TCQ 7'h00;
    trn_rerrfwd_prev   <= #TCQ 1'b0;
    trn_recrc_err_prev <= #TCQ 1'b0;
    trn_reof_prev      <= #TCQ 1'b0;
    trn_rsrc_dsc_prev  <= #TCQ 1'b0;
  end
  else begin
    // prev buffer works by checking trn_rdst_rdy. When trn_rdst_rdy is
    // asserted, a new value is present on the interface.
    if(trn_rdst_rdy) begin
      trn_rd_prev        <= #TCQ trn_rd_DW_swapped;
      trn_rsof_prev      <= #TCQ trn_rsof;
      trn_rrem_prev      <= #TCQ trn_rrem;
      trn_rbar_hit_prev  <= #TCQ trn_rbar_hit;
      trn_rerrfwd_prev   <= #TCQ trn_rerrfwd;
      trn_recrc_err_prev <= #TCQ trn_recrc_err;
      trn_rsrc_rdy_prev  <= #TCQ rsrc_rdy_filtered;
      trn_reof_prev      <= #TCQ trn_reof;
      trn_rsrc_dsc_prev  <= #TCQ trn_rsrc_dsc || dsc_flag;
    end
  end
end


//----------------------------------------------------------------------------//
// Create TDATA                                                               //
//----------------------------------------------------------------------------//

// Convert TRN data format to AXI data format. AXI is DWORD swapped from TRN
// 128-bit:                 64-bit:                  32-bit:
// TRN DW0 maps to AXI DW3  TRN DW0 maps to AXI DW1  TNR DW0 maps to AXI DW0
// TRN DW1 maps to AXI DW2  TRN DW1 maps to AXI DW0
// TRN DW2 maps to AXI DW1
// TRN DW3 maps to AXI DW0
generate
  if(C_DATA_WIDTH == 128) begin : rd_DW_swap_128
    assign trn_rd_DW_swapped = {trn_rd[31:0],
                                trn_rd[63:32],
                                trn_rd[95:64],
                                trn_rd[127:96]};
  end
  else if(C_DATA_WIDTH == 64) begin : rd_DW_swap_64
    assign trn_rd_DW_swapped = {trn_rd[31:0], trn_rd[63:32]};
  end
  else begin : rd_DW_swap_32
    assign trn_rd_DW_swapped = trn_rd;
  end
endgenerate


// Create special buffer which locks in the proper value of TDATA depending
// on whether the user is throttling or not. This buffer has three states:
//
//       HOLD state: TDATA maintains its current value
//                   - the user has throttled the PCIe block
//   PREVIOUS state: the buffer provides the previous value on trn_rd
//                   - the user has finished throttling, and is a little behind
//                     the PCIe block
//    CURRENT state: the buffer passes the current value on trn_rd
//                   - the user is caught up and ready to receive the latest
//                     data from the PCIe block
always @(posedge user_clk) begin
  if(user_rst) begin
    m_axis_rx_tdata <= #TCQ {C_DATA_WIDTH{1'b0}};
  end
  else begin
    if(!data_hold) begin
      // PREVIOUS state
      if(data_prev) begin
        m_axis_rx_tdata <= #TCQ trn_rd_prev;
      end

      // CURRENT state
      else begin
        m_axis_rx_tdata <= #TCQ trn_rd_DW_swapped;
      end
    end
    // else HOLD state
  end
end

// Logic to instruct pipeline to hold its value
assign data_hold = (!m_axis_rx_tready && m_axis_rx_tvalid);

// Logic to instruct pipeline to use previous bus values. Always use previous
// value after holding a value.
always @(posedge user_clk) begin
  if(user_rst) begin
    data_prev <= #TCQ 1'b0;
  end
  else begin
    data_prev <= #TCQ data_hold;
  end
end


//----------------------------------------------------------------------------//
// Create TVALID, TLAST, tkeep, TUSER                                         //
// -----------------------------------                                        //
// Use the same strategy for these signals as for TDATA, except here we need  //
// an extra provision for null packets.                                       //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    m_axis_rx_tvalid <= #TCQ 1'b0;
    reg_tlast        <= #TCQ 1'b0;
    reg_tkeep        <= #TCQ {KEEP_WIDTH{1'b1}};
    m_axis_rx_tuser  <= #TCQ 22'h0;
  end
  else begin
    if(!data_hold) begin
      // If in a null packet, use null generated value
      if(null_mux_sel) begin
        m_axis_rx_tvalid <= #TCQ null_rx_tvalid;
        reg_tlast        <= #TCQ null_rx_tlast;
        reg_tkeep        <= #TCQ null_rx_tkeep;
        m_axis_rx_tuser  <= #TCQ {null_is_eof, 17'h0000};
      end

      // PREVIOUS state
      else if(data_prev) begin
        m_axis_rx_tvalid <= #TCQ (trn_rsrc_rdy_prev || dsc_flag);
        reg_tlast        <= #TCQ trn_reof_prev;
        reg_tkeep        <= #TCQ tkeep_prev;
        m_axis_rx_tuser  <= #TCQ {is_eof_prev,          // TUSER bits [21:17]
                                  2'b00,                // TUSER bits [16:15]
                                  is_sof_prev,          // TUSER bits [14:10]
                                  1'b0,                 // TUSER bit  [9]
                                  trn_rbar_hit_prev,    // TUSER bits [8:2]
                                  trn_rerrfwd_prev,     // TUSER bit  [1]
                                  trn_recrc_err_prev};  // TUSER bit  [0]
      end

      // CURRENT state
      else begin
        m_axis_rx_tvalid <= #TCQ (rsrc_rdy_filtered || dsc_flag);
        reg_tlast        <= #TCQ trn_reof;
        reg_tkeep        <= #TCQ tkeep;
        m_axis_rx_tuser  <= #TCQ {is_eof,               // TUSER bits [21:17]
                                  2'b00,                // TUSER bits [16:15]
                                  is_sof,               // TUSER bits [14:10]
                                  1'b0,                 // TUSER bit  [9]
                                  trn_rbar_hit,         // TUSER bits [8:2]
                                  trn_rerrfwd,          // TUSER bit  [1]
                                  trn_recrc_err};       // TUSER bit  [0]
      end
    end
    // else HOLD state
  end
end

// Hook up TLAST and tkeep depending on interface width
generate
  // For 128-bit interface, don't pass TLAST and tkeep to user (is_eof and
  // is_data passed to user instead). reg_tlast is still used internally.
  if(C_DATA_WIDTH == 128) begin : tlast_tkeep_hookup_128
    assign m_axis_rx_tlast = 1'b0;
    assign m_axis_rx_tkeep = {KEEP_WIDTH{1'b1}};
  end

  // For 64/32-bit interface, pass TLAST to user.
  else begin : tlast_tkeep_hookup_64_32
    assign m_axis_rx_tlast = reg_tlast;
    assign m_axis_rx_tkeep = reg_tkeep;
  end
endgenerate


//----------------------------------------------------------------------------//
// Create tkeep                                                               //
// ------------                                                               //
// Convert RREM to STRB. Here, we are converting the encoding method for the  //
// location of the EOF from TRN flavor (rrem) to AXI (tkeep).                 //
//                                                                            //
// NOTE: for each configuration, we need two values of tkeep, the current and //
//       previous values. The need for these two values is described below.   //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : rrem_to_tkeep_128
    // TLAST and tkeep not used in 128-bit interface. is_sof and is_eof used
    // instead.
    assign tkeep      = 16'h0000;
    assign tkeep_prev = 16'h0000;
  end
  else if(C_DATA_WIDTH == 64) begin : rrem_to_tkeep_64
    // 64-bit interface: contains 2 DWORDs per cycle, for a total of 8 bytes
    //  - tkeep has only two possible values here, 0xFF or 0x0F
    assign tkeep      = trn_rrem      ? 8'hFF : 8'h0F;
    assign tkeep_prev = trn_rrem_prev ? 8'hFF : 8'h0F;
  end
  else begin : rrem_to_tkeep_32
    // 32-bit interface: contains 1 DWORD per cycle, for a total of 4 bytes
    //  - tkeep is always 0xF in this case, due to the nature of the PCIe block
    assign tkeep      = 4'hF;
    assign tkeep_prev = 4'hF;
  end
endgenerate


//----------------------------------------------------------------------------//
// Create is_sof                                                              //
// -------------                                                              //
// is_sof is a signal to the user indicating the location of SOF in TDATA   . //
// Due to inherent 64-bit alignment of packets from the block, the only       //
// possible values are:                                                       //
//                      Value                      Valid data widths          //
//                      5'b11000 (sof @ byte 8)    128                        //
//                      5'b10000 (sof @ byte 0)    128, 64, 32                //
//                      5'b00000 (sof not present) 128, 64, 32                //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : is_sof_128
    assign is_sof      = {(trn_rsof && !trn_rsrc_dsc), // bit 4:   enable
                          (trn_rsof && !trn_rrem[1]),  // bit 3:   sof @ byte 8?
                          3'b000};                     // bit 2-0: hardwired 0

    assign is_sof_prev = {(trn_rsof_prev && !trn_rsrc_dsc_prev), // bit 4
                          (trn_rsof_prev && !trn_rrem_prev[1]),  // bit 3
                          3'b000};                               // bit 2-0
  end
  else begin : is_sof_64_32
    assign is_sof      = {(trn_rsof && !trn_rsrc_dsc), // bit 4:   enable
                          4'b0000};                    // bit 3-0: hardwired 0

    assign is_sof_prev = {(trn_rsof_prev && !trn_rsrc_dsc_prev), // bit 4
                          4'b0000};                              // bit 3-0
  end
endgenerate


//----------------------------------------------------------------------------//
// Create is_eof                                                              //
// -------------                                                              //
// is_eof is a signal to the user indicating the location of EOF in TDATA   . //
// Due to DWORD granularity of packets from the block, the only               //
// possible values are:                                                       //
//                      Value                      Valid data widths          //
//                      5'b11111 (eof @ byte 15)   128                        //
//                      5'b11011 (eof @ byte 11)   128                        //
//                      5'b10111 (eof @ byte 7)    128, 64                    //
//                      5'b10011 (eof @ byte 3)`   128, 64, 32                //
//                      5'b00011 (eof not present) 128, 64, 32                //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : is_eof_128
    assign is_eof      = {trn_reof,      // bit 4:   enable
                          trn_rrem,      // bit 3-2: encoded eof loc rom block
                          2'b11};        // bit 1-0: hardwired 1

    assign is_eof_prev = {trn_reof_prev, // bit 4:   enable
                          trn_rrem_prev, // bit 3-2: encoded eof loc from block
                          2'b11};        // bit 1-0: hardwired 1
  end
  else if(C_DATA_WIDTH == 64) begin : is_eof_64
    assign is_eof      = {trn_reof,      // bit 4:   enable
                          1'b0,          // bit 3:   hardwired 0
                          trn_rrem,      // bit 2:   encoded eof loc from block
                          2'b11};        // bit 1-0: hardwired 1

    assign is_eof_prev = {trn_reof_prev, // bit 4:   enable
                          1'b0,          // bit 3:   hardwired 0
                          trn_rrem_prev, // bit 2:   encoded eof loc from block
                          2'b11};        // bit 1-0: hardwired 1
  end
  else begin : is_eof_32
    assign is_eof      = {trn_reof,      // bit 4:   enable
                          4'b0011};      // bit 3-0: hardwired to byte 3

    assign is_eof_prev = {trn_reof_prev, // bit 4:   enable
                          4'b0011};      // bit 3-0: hardwired to byte 3
  end
endgenerate



//----------------------------------------------------------------------------//
// Create trn_rdst_rdy                                                        //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    trn_rdst_rdy <= #TCQ 1'b0;
  end
  else begin
    // If in a null packet, use null generated value
    if(null_mux_sel && m_axis_rx_tready) begin
      trn_rdst_rdy <= #TCQ null_rdst_rdy;
    end

    // If a discontinue needs to be serviced, throttle the block until we are
    // ready to pad out the packet.
    else if(dsc_flag) begin
      trn_rdst_rdy <= #TCQ 1'b0;
    end

    // If in a packet, pass user back-pressure directly to block
    else if(m_axis_rx_tvalid) begin
      trn_rdst_rdy <= #TCQ m_axis_rx_tready;
    end

    // If idle, default to no back-pressure. We need to default to the
    // "ready to accept data" state to make sure we catch the first
    // clock of data of a new packet.
    else begin
      trn_rdst_rdy <= #TCQ 1'b1;
    end
  end
end

//----------------------------------------------------------------------------//
// Create null_mux_sel                                                        //
// null_mux_sel is the signal used to detect a discontinue situation and      //
// mux in the null packet generated in rx_null_gen. Only mux in null data     //
// when not at the beginningof a packet. SOF discontinues do not require      //
// padding, as the whole packet is simply squashed instead.                   //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    null_mux_sel <= #TCQ 1'b0;
  end
  else begin
    // NULL packet done
    if(null_mux_sel && null_rx_tlast && m_axis_rx_tready)
    begin
      null_mux_sel <= #TCQ 1'b0;
    end

    // Discontinue detected and we're in packet, so switch to NULL packet
    else if(dsc_flag && !data_hold) begin
      null_mux_sel <= #TCQ 1'b1;
    end
  end
end


//----------------------------------------------------------------------------//
// Create discontinue tracking signals                                        //
//----------------------------------------------------------------------------//
// Create signal trn_in_packet, which is needed to validate trn_rsrc_dsc. We
// should ignore trn_rsrc_dsc when it's asserted out-of-packet.
always @(posedge user_clk) begin
  if(user_rst) begin
    trn_in_packet <= #TCQ 1'b0;
  end
  else begin
    if(trn_rsof && !trn_reof && rsrc_rdy_filtered && trn_rdst_rdy)
    begin
      trn_in_packet <= #TCQ 1'b1;
    end
    else if(trn_rsrc_dsc) begin
      trn_in_packet <= #TCQ 1'b0;
    end
    else if(trn_reof && !trn_rsof && trn_rsrc_rdy && trn_rdst_rdy) begin
      trn_in_packet <= #TCQ 1'b0;
    end
  end
end


// Create dsc_flag, which identifies and stores mid-packet discontinues that
// require null packet padding. This signal is edge sensitive to trn_rsrc_dsc,
// to make sure we don't service the same dsc twice in the event that
// trn_rsrc_dsc stays asserted for longer than it takes to pad out the packet.
assign dsc_detect = trn_rsrc_dsc && !trn_rsrc_dsc_d && trn_in_packet &&
                         (!trn_rsof || trn_reof) && !(trn_rdst_rdy && trn_reof);

always @(posedge user_clk) begin
  if(user_rst) begin
    reg_dsc_detect <= #TCQ 1'b0;
    trn_rsrc_dsc_d <= #TCQ 1'b0;
  end
  else begin
    if(dsc_detect) begin
      reg_dsc_detect <= #TCQ 1'b1;
    end
    else if(null_mux_sel) begin
      reg_dsc_detect <= #TCQ 1'b0;
    end

    trn_rsrc_dsc_d <= #TCQ trn_rsrc_dsc;
  end
end

assign dsc_flag = dsc_detect || reg_dsc_detect;



//----------------------------------------------------------------------------//
// Create np_counter (V6 128-bit only). This counter tells the V6 128-bit     //
// interface core how many NP packets have left the RX pipeline. The V6       //
// 128-bit interface uses this count to perform rnp_ok modulation.            //
//----------------------------------------------------------------------------//
generate
  if(C_FAMILY == "V6" && C_DATA_WIDTH == 128) begin : np_cntr_to_128_enabled
    reg [2:0] reg_np_counter;

    // Look for NP packets beginning on lower (i.e. unaligned) start
    wire mrd_lower      = (!(|m_axis_rx_tdata[92:88]) && !m_axis_rx_tdata[94]);
    wire mrd_lk_lower   = (m_axis_rx_tdata[92:88] == 5'b00001);
    wire io_rdwr_lower  = (m_axis_rx_tdata[92:88] == 5'b00010);
    wire cfg_rdwr_lower = (m_axis_rx_tdata[92:89] == 4'b0010);
    wire atomic_lower   = ((&m_axis_rx_tdata[91:90]) && m_axis_rx_tdata[94]);

    wire np_pkt_lower = (mrd_lower      ||
                         mrd_lk_lower   ||
                         io_rdwr_lower  ||
                         cfg_rdwr_lower ||
                         atomic_lower) && m_axis_rx_tuser[13];

    // Look for NP packets beginning on upper (i.e. aligned) start
    wire mrd_upper      = (!(|m_axis_rx_tdata[28:24]) && !m_axis_rx_tdata[30]);
    wire mrd_lk_upper   = (m_axis_rx_tdata[28:24] == 5'b00001);
    wire io_rdwr_upper  = (m_axis_rx_tdata[28:24] == 5'b00010);
    wire cfg_rdwr_upper = (m_axis_rx_tdata[28:25] == 4'b0010);
    wire atomic_upper   = ((&m_axis_rx_tdata[27:26]) && m_axis_rx_tdata[30]);

    wire np_pkt_upper = (mrd_upper      ||
                         mrd_lk_upper   ||
                         io_rdwr_upper  ||
                         cfg_rdwr_upper ||
                         atomic_upper) && !m_axis_rx_tuser[13];

    wire pkt_accepted =
                    m_axis_rx_tuser[14] && m_axis_rx_tready && m_axis_rx_tvalid;

    // Increment counter whenever an NP packet leaves the RX pipeline
    always @(posedge user_clk)  begin
      if (user_rst) begin
        reg_np_counter <= #TCQ 0;
      end
      else begin
        if((np_pkt_lower || np_pkt_upper) && pkt_accepted)
        begin
          reg_np_counter <= #TCQ reg_np_counter + 3'h1;
        end
      end
    end

    assign np_counter = reg_np_counter;
  end
  else begin : np_cntr_to_128_disabled
    assign np_counter = 3'h0;
  end
endgenerate


endmodule



`timescale 1ns/1ps
module model_ap2_tst_axi_basic_rx_null_gen # (
  parameter C_DATA_WIDTH = 128,           // RX/TX interface data width
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8            // KEEP width
  ) (

  // AXI RX
  //-----------
  input      [C_DATA_WIDTH-1:0] m_axis_rx_tdata,     // RX data to user
  input                         m_axis_rx_tvalid,    // RX data is valid
  input                         m_axis_rx_tready,    // RX ready for data
  input                         m_axis_rx_tlast,     // RX data is last
  input                  [21:0] m_axis_rx_tuser,     // RX user signals

  // Null Inputs
  //-----------
  output                        null_rx_tvalid,      // NULL generated tvalid
  output                        null_rx_tlast,       // NULL generated tlast
  output       [KEEP_WIDTH-1:0] null_rx_tkeep,       // NULL generated tkeep
  output                        null_rdst_rdy,       // NULL generated rdst_rdy
  output reg              [4:0] null_is_eof,         // NULL generated is_eof

  // System
  //-----------
  input                         user_clk,            // user clock from block
  input                         user_rst             // user reset from block
);


localparam INTERFACE_WIDTH_DWORDS = (C_DATA_WIDTH == 128) ? 11'd4 :
                                           (C_DATA_WIDTH == 64) ? 11'd2 : 11'd1;

//----------------------------------------------------------------------------//
// NULL packet generator state machine                                        //
// This state machine shadows the AXI RX interface, tracking each packet as   //
// it's passed to the AXI user. When a multi-cycle packet is detected, the    //
// state machine automatically generates a "null" packet. In the event of a   //
// discontinue, the RX pipeline can switch over to this null packet as        //
// necessary.                                                                 //
//----------------------------------------------------------------------------//

// State machine variables and states
localparam            IDLE      = 0;
localparam            IN_PACKET = 1;
reg                   cur_state;
reg                   next_state;

// Signals for tracking a packet on the AXI interface
reg            [11:0] reg_pkt_len_counter;
reg            [11:0] pkt_len_counter;
wire           [11:0] pkt_len_counter_dec;
wire                  pkt_done;

// Calculate packet fields, which are needed to determine total packet length.
wire           [11:0] new_pkt_len;
wire            [9:0] payload_len;
wire            [1:0] packet_fmt;
wire                  packet_td;
reg             [3:0] packet_overhead;

// Misc.
wire [KEEP_WIDTH-1:0] eof_tkeep;
wire                  straddle_sof;
wire                  eof;


// Create signals to detect sof and eof situations. These signals vary depending
// on data width.
assign eof = m_axis_rx_tuser[21];
generate
  if(C_DATA_WIDTH == 128) begin : sof_eof_128
    assign straddle_sof = (m_axis_rx_tuser[14:13] == 2'b11);
  end
  else begin : sof_eof_64_32
    assign straddle_sof = 1'b0;
  end
endgenerate


//----------------------------------------------------------------------------//
// Calculate the length of the packet being presented on the RX interface. To //
// do so, we need the relevent packet fields that impact total packet length. //
// These are:                                                                 //
//   - Header length: obtained from bit 1 of FMT field in 1st DWORD of header //
//   - Payload length: obtained from LENGTH field in 1st DWORD of header      //
//   - TLP digest: obtained from TD field in 1st DWORD of header              //
//   - Current data: the number of bytes that have already been presented     //
//                   on the data interface                                    //
//                                                                            //
// packet length = header + payload + tlp digest - # of DWORDS already        //
//                 transmitted                                                //
//                                                                            //
// packet_overhead is where we calculate everything except payload.           //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : len_calc_128
    assign packet_fmt  = straddle_sof ?
                                m_axis_rx_tdata[94:93] : m_axis_rx_tdata[30:29];
    assign packet_td   = straddle_sof ?
                                      m_axis_rx_tdata[79] : m_axis_rx_tdata[15];
    assign payload_len = packet_fmt[1] ?
         (straddle_sof ? m_axis_rx_tdata[73:64] : m_axis_rx_tdata[9:0]) : 10'h0;

    always @(*) begin
      // In 128-bit mode, the amount of data currently on the interface
      // depends on whether we're straddling or not. If so, 2 DWORDs have been
      // seen. If not, 4 DWORDs.
      case({packet_fmt[0], packet_td, straddle_sof})
        //                        Header +  TD  - Data currently on interface
        3'b0_0_0: packet_overhead = 4'd3 + 4'd0 - 4'd4;
        3'b0_0_1: packet_overhead = 4'd3 + 4'd0 - 4'd2;
        3'b0_1_0: packet_overhead = 4'd3 + 4'd1 - 4'd4;
        3'b0_1_1: packet_overhead = 4'd3 + 4'd1 - 4'd2;
        3'b1_0_0: packet_overhead = 4'd4 + 4'd0 - 4'd4;
        3'b1_0_1: packet_overhead = 4'd4 + 4'd0 - 4'd2;
        3'b1_1_0: packet_overhead = 4'd4 + 4'd1 - 4'd4;
        3'b1_1_1: packet_overhead = 4'd4 + 4'd1 - 4'd2;
      endcase
    end
assign new_pkt_len =
         {{9{packet_overhead[3]}}, packet_overhead[2:0]} + {2'b0, payload_len};
  end
  else if(C_DATA_WIDTH == 64) begin : len_calc_64
    assign packet_fmt  = m_axis_rx_tdata[30:29];
    assign packet_td   = m_axis_rx_tdata[15];
    assign payload_len = packet_fmt[1] ? m_axis_rx_tdata[9:0] : 10'h0;

    always @(*) begin
      // 64-bit mode: no straddling, so always 2 DWORDs
      case({packet_fmt[0], packet_td})
        //                      Header +  TD  - Data currently on interface
        2'b0_0: packet_overhead[1:0] = 2'b01 ;//4'd3 + 4'd0 - 4'd2; // 1
        2'b0_1: packet_overhead[1:0] = 2'b10 ;//4'd3 + 4'd1 - 4'd2; // 2
        2'b1_0: packet_overhead[1:0] = 2'b10 ;//4'd4 + 4'd0 - 4'd2; // 2 
        2'b1_1: packet_overhead[1:0] = 2'b11 ;//4'd4 + 4'd1 - 4'd2; // 3
      endcase
    end
assign new_pkt_len =
         {{10{1'b0}}, packet_overhead[1:0]} + {2'b0, payload_len};
  end
  else begin : len_calc_32
    assign packet_fmt  = m_axis_rx_tdata[30:29];
    assign packet_td   = m_axis_rx_tdata[15];
    assign payload_len = packet_fmt[1] ? m_axis_rx_tdata[9:0] : 10'h0;

    always @(*) begin
      // 32-bit mode: no straddling, so always 1 DWORD
      case({packet_fmt[0], packet_td})
        //                      Header +  TD  - Data currently on interface
        2'b0_0: packet_overhead = 4'd3 + 4'd0 - 4'd1;
        2'b0_1: packet_overhead = 4'd3 + 4'd1 - 4'd1;
        2'b1_0: packet_overhead = 4'd4 + 4'd0 - 4'd1;
        2'b1_1: packet_overhead = 4'd4 + 4'd1 - 4'd1;
      endcase
    end
assign new_pkt_len =
         {{9{packet_overhead[3]}}, packet_overhead[2:0]} + {2'b0, payload_len};
  end
endgenerate

// Now calculate actual packet length, adding the packet overhead and the
// payload length. This is signed math, so sign-extend packet_overhead.
// NOTE: a payload length of zero means 1024 DW in the PCIe spec, but this
//       behavior isn't supported in our block.
//assign new_pkt_len =
//         {{9{packet_overhead[3]}}, packet_overhead[2:0]} + {2'b0, payload_len};


// Math signals needed in the state machine below. These are seperate wires to
// help ensure synthesis tools sre smart about optimizing them.
assign pkt_len_counter_dec = reg_pkt_len_counter - INTERFACE_WIDTH_DWORDS;
assign pkt_done = (reg_pkt_len_counter <= INTERFACE_WIDTH_DWORDS);

//----------------------------------------------------------------------------//
// Null generator Mealy state machine. Determine outputs based on:            //
//   1) current st                                                            //
//   2) current inp                                                           //
//----------------------------------------------------------------------------//
always @(*) begin
  case (cur_state)

    // IDLE state: the interface is IDLE and we're waiting for a packet to
    // start. If a packet starts, move to state IN_PACKET and begin tracking
    // it as long as it's NOT a single cycle packet (indicated by assertion of
    // eof at packet start)
    IDLE: begin
      if(m_axis_rx_tvalid && m_axis_rx_tready && !eof) begin
        next_state = IN_PACKET;
      end
      else begin
        next_state = IDLE;
      end

      pkt_len_counter = new_pkt_len;
    end

    // IN_PACKET: a mutli-cycle packet is in progress and we're tracking it. We
    // are in lock-step with the AXI interface decrementing our packet length
    // tracking reg, and waiting for the packet to finish.
    //
    // * If packet finished and a new one starts, this is a straddle situation.
    //   Next state is IN_PACKET (128-bit only).
    // * If the current packet is done, next state is IDLE.
    // * Otherwise, next state is IN_PACKET.
    IN_PACKET: begin
      // Straddle packet
      if((C_DATA_WIDTH == 128) && straddle_sof && m_axis_rx_tvalid) begin
        pkt_len_counter = new_pkt_len;
        next_state = IN_PACKET;
      end

      // Current packet finished
      else if(m_axis_rx_tready && pkt_done)
      begin
        pkt_len_counter = new_pkt_len;
        next_state      = IDLE;
      end

      // Packet in progress
      else begin
        if(m_axis_rx_tready) begin
          // Not throttled
          pkt_len_counter = pkt_len_counter_dec;
        end
        else begin
          // Throttled
          pkt_len_counter = reg_pkt_len_counter;
        end

        next_state = IN_PACKET;
      end
    end

    default: begin
      pkt_len_counter = reg_pkt_len_counter;
      next_state      = IDLE;
    end
  endcase
end


// Synchronous NULL packet generator state machine logic
always @(posedge user_clk) begin
  if(user_rst) begin
    cur_state           <= #TCQ IDLE;
    reg_pkt_len_counter <= #TCQ 12'h0;
  end
  else begin
    cur_state           <= #TCQ next_state;
    reg_pkt_len_counter <= #TCQ pkt_len_counter;
  end
end


// Generate tkeep/is_eof for an end-of-packet situation.
generate
  if(C_DATA_WIDTH == 128) begin : strb_calc_128
    always @(*) begin
      // Assign null_is_eof depending on how many DWORDs are left in the
      // packet.
      case(pkt_len_counter)
        10'd1:   null_is_eof = 5'b10011;
        10'd2:   null_is_eof = 5'b10111;
        10'd3:   null_is_eof = 5'b11011;
        10'd4:   null_is_eof = 5'b11111;
        default: null_is_eof = 5'b00011;
      endcase
    end

    // tkeep not used in 128-bit interface
    assign eof_tkeep = {KEEP_WIDTH{1'b0}};
  end
  else if(C_DATA_WIDTH == 64) begin : strb_calc_64
    always @(*) begin
      // Assign null_is_eof depending on how many DWORDs are left in the
      // packet.
      case(pkt_len_counter)
        10'd1:   null_is_eof = 5'b10011;
        10'd2:   null_is_eof = 5'b10111;
        default: null_is_eof = 5'b00011;
      endcase
    end

    // Assign tkeep to 0xFF or 0x0F depending on how many DWORDs are left in
    // the current packet.
    assign eof_tkeep = { ((pkt_len_counter == 12'd2) ? 4'hF:4'h0), 4'hF };
  end
  else begin : strb_calc_32
    always @(*) begin
      // is_eof is either on or off for 32-bit
      if(pkt_len_counter == 12'd1) begin
        null_is_eof = 5'b10011;
      end
      else begin
        null_is_eof = 5'b00011;
      end
    end

    // The entire DWORD is always valid in 32-bit mode, so tkeep is always 0xF
    assign eof_tkeep = 4'hF;
  end
endgenerate


// Finally, use everything we've generated to calculate our NULL outputs
assign null_rx_tvalid = 1'b1;
assign null_rx_tlast  = (pkt_len_counter <= INTERFACE_WIDTH_DWORDS);
assign null_rx_tkeep  = null_rx_tlast ? eof_tkeep : {KEEP_WIDTH{1'b1}};
assign null_rdst_rdy  = null_rx_tlast;

endmodule


`timescale 1ns/1ps
module model_ap2_tst_axi_basic_tx #(
  parameter C_DATA_WIDTH  = 128,          // RX/TX interface data width
  parameter C_FAMILY      = "X7",         // Targeted FPGA family
  parameter C_ROOT_PORT   = "FALSE",      // PCIe block is in root port mode
  parameter C_PM_PRIORITY = "FALSE",      // Disable TX packet boundary thrtl
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter REM_WIDTH  = (C_DATA_WIDTH == 128) ? 2 : 1, // trem/rrem width
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8               // KEEP width
  ) (
  //---------------------------------------------//
  // User Design I/O                             //
  //---------------------------------------------//

  // AXI TX
  //-----------
  input   [C_DATA_WIDTH-1:0] s_axis_tx_tdata,        // TX data from user
  input                      s_axis_tx_tvalid,       // TX data is valid
  output                     s_axis_tx_tready,       // TX ready for data
  input     [KEEP_WIDTH-1:0] s_axis_tx_tkeep,        // TX strobe byte enables
  input                      s_axis_tx_tlast,        // TX data is last
  input                [3:0] s_axis_tx_tuser,        // TX user signals

  // User Misc.
  //-----------
  input                      user_turnoff_ok,        // Turnoff OK from user
  input                      user_tcfg_gnt,          // Send cfg OK from user

  //---------------------------------------------//
  // PCIe Block I/O                              //
  //---------------------------------------------//

  // TRN TX
  //-----------
  output [C_DATA_WIDTH-1:0] trn_td,                  // TX data from block
  output                    trn_tsof,                // TX start of packet
  output                    trn_teof,                // TX end of packet
  output                    trn_tsrc_rdy,            // TX source ready
  input                     trn_tdst_rdy,            // TX destination ready
  output                    trn_tsrc_dsc,            // TX source discontinue
  output    [REM_WIDTH-1:0] trn_trem,                // TX remainder
  output                    trn_terrfwd,             // TX error forward
  output                    trn_tstr,                // TX streaming enable
  input               [5:0] trn_tbuf_av,             // TX buffers available
  output                    trn_tecrc_gen,           // TX ECRC generate

  // TRN Misc.
  //-----------
  input                     trn_tcfg_req,            // TX config request
  output                    trn_tcfg_gnt,            // RX config grant
  input                     trn_lnk_up,              // PCIe link up

  // 7 Series/Virtex6 PM
  //-----------
  input               [2:0] cfg_pcie_link_state,     // Encoded PCIe link state

  // Virtex6 PM
  //-----------
  input                     cfg_pm_send_pme_to,      // PM send PME turnoff msg
  input               [1:0] cfg_pmcsr_powerstate,    // PMCSR power state
  input              [31:0] trn_rdllp_data,          // RX DLLP data
  input                     trn_rdllp_src_rdy,       // RX DLLP source ready

  // Virtex6/Spartan6 PM
  //-----------
  input                     cfg_to_turnoff,          // Turnoff request
  output                    cfg_turnoff_ok,          // Turnoff grant

  // System
  //-----------
  input                     user_clk,                // user clock from block
  input                     user_rst                 // user reset from block
);


wire tready_thrtl;

//---------------------------------------------//
// TX Data Pipeline                            //
//---------------------------------------------//

model_ap2_tst_axi_basic_tx_pipeline #(
  .C_DATA_WIDTH( C_DATA_WIDTH ),
  .C_PM_PRIORITY( C_PM_PRIORITY ),
  .TCQ( TCQ ),

  .REM_WIDTH( REM_WIDTH ),
  .KEEP_WIDTH( KEEP_WIDTH )
) model_ap2_tst_tx_pipeline_inst (

  // Incoming AXI RX
  //-----------
  .s_axis_tx_tdata( s_axis_tx_tdata ),
  .s_axis_tx_tready( s_axis_tx_tready ),
  .s_axis_tx_tvalid( s_axis_tx_tvalid ),
  .s_axis_tx_tkeep( s_axis_tx_tkeep ),
  .s_axis_tx_tlast( s_axis_tx_tlast ),
  .s_axis_tx_tuser( s_axis_tx_tuser ),

  // Outgoing TRN TX
  //-----------
  .trn_td( trn_td ),
  .trn_tsof( trn_tsof ),
  .trn_teof( trn_teof ),
  .trn_tsrc_rdy( trn_tsrc_rdy ),
  .trn_tdst_rdy( trn_tdst_rdy ),
  .trn_tsrc_dsc( trn_tsrc_dsc ),
  .trn_trem( trn_trem ),
  .trn_terrfwd( trn_terrfwd ),
  .trn_tstr( trn_tstr ),
  .trn_tecrc_gen( trn_tecrc_gen ),
  .trn_lnk_up( trn_lnk_up ),

  // System
  //-----------
  .tready_thrtl( tready_thrtl ),
  .user_clk( user_clk ),
  .user_rst( user_rst )
);


//---------------------------------------------//
// TX Throttle Controller                      //
//---------------------------------------------//

generate
  if(C_PM_PRIORITY == "FALSE") begin : thrtl_ctl_enabled
model_ap2_tst_axi_basic_tx_thrtl_ctl #(
      .C_DATA_WIDTH( C_DATA_WIDTH ),
      .C_FAMILY( C_FAMILY ),
      .C_ROOT_PORT( C_ROOT_PORT ),
      .TCQ( TCQ )

    ) model_ap2_tst_tx_thrl_ctl_inst (

      // Outgoing AXI TX
      //-----------
      .s_axis_tx_tdata( s_axis_tx_tdata ),
      .s_axis_tx_tvalid( s_axis_tx_tvalid ),
      .s_axis_tx_tuser( s_axis_tx_tuser ),
      .s_axis_tx_tlast( s_axis_tx_tlast ),

      // User Misc.
      //-----------
      .user_turnoff_ok( user_turnoff_ok ),
      .user_tcfg_gnt( user_tcfg_gnt ),

      // Incoming TRN RX
      //-----------
      .trn_tbuf_av( trn_tbuf_av ),
      .trn_tdst_rdy( trn_tdst_rdy ),

      // TRN Misc.
      //-----------
      .trn_tcfg_req( trn_tcfg_req ),
      .trn_tcfg_gnt( trn_tcfg_gnt ),
      .trn_lnk_up( trn_lnk_up ),

      // 7 Seriesq/Virtex6 PM
      //-----------
      .cfg_pcie_link_state( cfg_pcie_link_state ),

      // Virtex6 PM
      //-----------
      .cfg_pm_send_pme_to( cfg_pm_send_pme_to ),
      .cfg_pmcsr_powerstate( cfg_pmcsr_powerstate ),
      .trn_rdllp_data( trn_rdllp_data ),
      .trn_rdllp_src_rdy( trn_rdllp_src_rdy ),

      // Spartan6 PM
      //-----------
      .cfg_to_turnoff( cfg_to_turnoff ),
      .cfg_turnoff_ok( cfg_turnoff_ok ),

      // System
      //-----------
      .tready_thrtl( tready_thrtl ),
      .user_clk( user_clk ),
      .user_rst( user_rst )
    );
  end
  else begin : thrtl_ctl_disabled
    assign tready_thrtl   = 1'b0;

    assign cfg_turnoff_ok = user_turnoff_ok;
    assign trn_tcfg_gnt   = user_tcfg_gnt;
  end
endgenerate

endmodule



`timescale 1ns/1ps
module model_ap2_tst_axi_basic_tx_pipeline #(
  parameter C_DATA_WIDTH = 128,           // RX/TX interface data width
  parameter C_PM_PRIORITY = "FALSE",      // Disable TX packet boundary thrtl
  parameter TCQ = 1,                      // Clock to Q time

  // Do not override parameters below this line
  parameter REM_WIDTH  = (C_DATA_WIDTH == 128) ? 2 : 1, // trem/rrem width
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8               // KEEP width
  ) (
  //---------------------------------------------//
  // User Design I/O                             //
  //---------------------------------------------//

  // AXI TX
  //-----------
  input      [C_DATA_WIDTH-1:0] s_axis_tx_tdata,     // TX data from user
  input                         s_axis_tx_tvalid,    // TX data is valid
  output                        s_axis_tx_tready,    // TX ready for data
  input        [KEEP_WIDTH-1:0] s_axis_tx_tkeep,     // TX strobe byte enables
  input                         s_axis_tx_tlast,     // TX data is last
  input                   [3:0] s_axis_tx_tuser,     // TX user signals

  //---------------------------------------------//
  // PCIe Block I/O                              //
  //---------------------------------------------//

  // TRN TX
  //-----------
  output     [C_DATA_WIDTH-1:0] trn_td,              // TX data from block
  output                        trn_tsof,            // TX start of packet
  output                        trn_teof,            // TX end of packet
  output                        trn_tsrc_rdy,        // TX source ready
  input                         trn_tdst_rdy,        // TX destination ready
  output                        trn_tsrc_dsc,        // TX source discontinue
  output        [REM_WIDTH-1:0] trn_trem,            // TX remainder
  output                        trn_terrfwd,         // TX error forward
  output                        trn_tstr,            // TX streaming enable
  output                        trn_tecrc_gen,       // TX ECRC generate
  input                         trn_lnk_up,          // PCIe link up

  // System
  //-----------
  input                         tready_thrtl,        // TREADY from thrtl ctl
  input                         user_clk,            // user clock from block
  input                         user_rst             // user reset from block
);


// Input register stage
reg  [C_DATA_WIDTH-1:0] reg_tdata;
reg                     reg_tvalid;
reg    [KEEP_WIDTH-1:0] reg_tkeep;
reg               [3:0] reg_tuser;
reg                     reg_tlast;
reg                     reg_tready;

// Pipeline utility signals
reg                     trn_in_packet;
reg                     axi_in_packet;
reg                     flush_axi;
wire                    disable_trn;
reg                     reg_disable_trn;

wire                    axi_beat_live  = s_axis_tx_tvalid && s_axis_tx_tready;
wire                    axi_end_packet = axi_beat_live && s_axis_tx_tlast;


//----------------------------------------------------------------------------//
// Convert TRN data format to AXI data format. AXI is DWORD swapped from TRN. //
// 128-bit:                 64-bit:                  32-bit:                  //
// TRN DW0 maps to AXI DW3  TRN DW0 maps to AXI DW1  TNR DW0 maps to AXI DW0  //
// TRN DW1 maps to AXI DW2  TRN DW1 maps to AXI DW0                           //
// TRN DW2 maps to AXI DW1                                                    //
// TRN DW3 maps to AXI DW0                                                    //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : td_DW_swap_128
    assign trn_td = {reg_tdata[31:0],
                     reg_tdata[63:32],
                     reg_tdata[95:64],
                     reg_tdata[127:96]};
  end
  else if(C_DATA_WIDTH == 64) begin : td_DW_swap_64
    assign trn_td = {reg_tdata[31:0], reg_tdata[63:32]};
  end
  else begin : td_DW_swap_32
    assign trn_td = reg_tdata;
  end
endgenerate


//----------------------------------------------------------------------------//
// Create trn_tsof. If we're not currently in a packet and TVALID goes high,  //
// assert TSOF.                                                               //
//----------------------------------------------------------------------------//
assign trn_tsof = reg_tvalid && !trn_in_packet;


//----------------------------------------------------------------------------//
// Create trn_in_packet. This signal tracks if the TRN interface is currently //
// in the middle of a packet, which is needed to generate trn_tsof            //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    trn_in_packet <= #TCQ 1'b0;
  end
  else begin
    if(trn_tsof && trn_tsrc_rdy && trn_tdst_rdy && !trn_teof) begin
      trn_in_packet <= #TCQ 1'b1;
    end
    else if((trn_in_packet && trn_teof && trn_tsrc_rdy) || !trn_lnk_up) begin
      trn_in_packet <= #TCQ 1'b0;
    end
  end
end


//----------------------------------------------------------------------------//
// Create axi_in_packet. This signal tracks if the AXI interface is currently //
// in the middle of a packet, which is needed in case the link goes down.     //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    axi_in_packet <= #TCQ 1'b0;
  end
  else begin
    if(axi_beat_live && !s_axis_tx_tlast) begin
      axi_in_packet <= #TCQ 1'b1;
    end
    else if(axi_beat_live) begin
      axi_in_packet <= #TCQ 1'b0;
    end
  end
end


//----------------------------------------------------------------------------//
// Create disable_trn. This signal asserts when the link goes down and        //
// triggers the deassertiong of trn_tsrc_rdy. The deassertion of disable_trn  //
// depends on C_PM_PRIORITY, as described below.                              //
//----------------------------------------------------------------------------//
generate
  // In the C_PM_PRIORITY pipeline, we disable the TRN interfacefrom the time
  // the link goes down until the the AXI interface is ready to accept packets
  // again (via assertion of TREADY). By waiting for TREADY, we allow the
  // previous value buffer to fill, so we're ready for any throttling by the
  // user or the block.
  if(C_PM_PRIORITY == "TRUE") begin : pm_priority_trn_flush
    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_disable_trn    <= #TCQ 1'b1;
      end
      else begin
        // When the link goes down, disable the TRN interface.
        if(!trn_lnk_up)
        begin
          reg_disable_trn  <= #TCQ 1'b1;
        end

        // When the link comes back up and the AXI interface is ready, we can
        // release the pipeline and return to normal operation.
        else if(!flush_axi && s_axis_tx_tready) begin
          reg_disable_trn <= #TCQ 1'b0;
        end
      end
    end

    assign disable_trn = reg_disable_trn;
  end

  // In the throttle-controlled pipeline, we don't have a previous value buffer.
  // The throttle control mechanism handles TREADY, so all we need to do is
  // detect when the link goes down and disable the TRN interface until the link
  // comes back up and the AXI interface is finished flushing any packets.
  else begin : thrtl_ctl_trn_flush
    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_disable_trn    <= #TCQ 1'b0;
      end
      else begin
        // If the link is down and AXI is in packet, disable TRN and look for
        // the end of the packet
        if(axi_in_packet && !trn_lnk_up && !axi_end_packet)
        begin
          reg_disable_trn  <= #TCQ 1'b1;
        end

        // AXI packet is ending, so we're done flushing
        else if(axi_end_packet) begin
          reg_disable_trn <= #TCQ 1'b0;
        end
      end
    end

    // Disable the TRN interface if link is down or we're still flushing the AXI
    // interface.
    assign disable_trn = reg_disable_trn || !trn_lnk_up;
  end
endgenerate


//----------------------------------------------------------------------------//
// Convert STRB to RREM. Here, we are converting the encoding method for the  //
// location of the EOF from AXI (tkeep) to TRN flavor (rrem).                 //
//----------------------------------------------------------------------------//
generate
  if(C_DATA_WIDTH == 128) begin : tkeep_to_trem_128
    //---------------------------------------//
    // Conversion table:                     //
    // trem    | tkeep                       //
    // [1] [0] | [15:12] [11:8] [7:4] [3:0]  //
    // ------------------------------------- //
    //  1   1  |   D3      D2    D1    D0    //
    //  1   0  |   --      D2    D1    D0    //
    //  0   1  |   --      --    D1    D0    //
    //  0   0  |   --      --    --    D0    //
    //---------------------------------------//

    wire   axi_DW_1    = reg_tkeep[7];
    wire   axi_DW_2    = reg_tkeep[11];
    wire   axi_DW_3    = reg_tkeep[15];
    assign trn_trem[1] = axi_DW_2;
    assign trn_trem[0] = axi_DW_3 || (axi_DW_1 && !axi_DW_2);
  end
  else if(C_DATA_WIDTH == 64) begin : tkeep_to_trem_64
    assign trn_trem    = reg_tkeep[7];
  end
  else begin : tkeep_to_trem_32
    assign trn_trem    = 1'b0;
  end
endgenerate


//----------------------------------------------------------------------------//
// Create remaining TRN signals                                               //
//----------------------------------------------------------------------------//
assign trn_teof      = reg_tlast;
assign trn_tecrc_gen = reg_tuser[0];
assign trn_terrfwd   = reg_tuser[1];
assign trn_tstr      = reg_tuser[2];
assign trn_tsrc_dsc  = reg_tuser[3];


//----------------------------------------------------------------------------//
// Pipeline stage                                                             //
//----------------------------------------------------------------------------//
// We need one of two approaches for the pipeline stage depending on the
// C_PM_PRIORITY parameter.
generate
  reg reg_tsrc_rdy;

  // If set to FALSE, that means the user wants to use the TX packet boundary
  // throttling feature. Since all Block throttling will now be predicted, we
  // can use a simple straight-through pipeline.
  if(C_PM_PRIORITY == "FALSE") begin : throttle_ctl_pipeline
    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_tdata        <= #TCQ {C_DATA_WIDTH{1'b0}};
        reg_tvalid       <= #TCQ 1'b0;
        reg_tkeep        <= #TCQ {KEEP_WIDTH{1'b0}};
        reg_tlast        <= #TCQ 1'b0;
        reg_tuser        <= #TCQ 4'h0;
        reg_tsrc_rdy     <= #TCQ 1'b0;
      end
      else begin
        reg_tdata        <= #TCQ s_axis_tx_tdata;
        reg_tvalid       <= #TCQ s_axis_tx_tvalid;
        reg_tkeep        <= #TCQ s_axis_tx_tkeep;
        reg_tlast        <= #TCQ s_axis_tx_tlast;
        reg_tuser        <= #TCQ s_axis_tx_tuser;

        // Hold trn_tsrc_rdy low when flushing a packet.
        reg_tsrc_rdy     <= #TCQ axi_beat_live && !disable_trn;
      end
    end

    assign trn_tsrc_rdy = reg_tsrc_rdy;

    // With TX packet boundary throttling, TREADY is pipelined in
    // axi_basic_tx_thrtl_ctl and wired through here.
    assign s_axis_tx_tready = tready_thrtl;
  end

  //**************************************************************************//

  // If C_PM_PRIORITY is set to TRUE, that means the user prefers to have all PM
  // functionality intact isntead of TX packet boundary throttling. Now the
  // Block could back-pressure at any time, which creates the standard problem
  // of potential data loss due to the handshaking latency. Here we need a
  // previous value buffer, just like the RX data path.
  else begin : pm_prioity_pipeline
    reg  [C_DATA_WIDTH-1:0] tdata_prev;
    reg                     tvalid_prev;
    reg    [KEEP_WIDTH-1:0] tkeep_prev;
    reg                     tlast_prev;
    reg               [3:0] tuser_prev;
    reg                     reg_tdst_rdy;

    wire                    data_hold;
    reg                     data_prev;


    //------------------------------------------------------------------------//
    // Previous value buffer                                                  //
    // ---------------------                                                  //
    // We are inserting a pipeline stage in between AXI and TRN, which causes //
    // some issues with handshaking signals trn_tsrc_rdy/s_axis_tx_tready.    //
    // The added cycle of latency in the path causes the Block to fall behind //
    // the AXI interface whenever it throttles.                               //
    //                                                                        //
    // To avoid loss of data, we must keep the previous value of all          //
    // s_axis_tx_* signals in case the Block throttles.                       //
    //------------------------------------------------------------------------//
    always @(posedge user_clk) begin
      if(user_rst) begin
        tdata_prev   <= #TCQ {C_DATA_WIDTH{1'b0}};
        tvalid_prev  <= #TCQ 1'b0;
        tkeep_prev   <= #TCQ {KEEP_WIDTH{1'b0}};
        tlast_prev   <= #TCQ 1'b0;
        tuser_prev   <= #TCQ 4'h 0;
      end
      else begin
        // prev buffer works by checking s_axis_tx_tready. When
        // s_axis_tx_tready is asserted, a new value is present on the
        // interface.
        if(!s_axis_tx_tready) begin
          tdata_prev   <= #TCQ tdata_prev;
          tvalid_prev  <= #TCQ tvalid_prev;
          tkeep_prev   <= #TCQ tkeep_prev;
          tlast_prev   <= #TCQ tlast_prev;
          tuser_prev   <= #TCQ tuser_prev;
        end
        else begin
          tdata_prev   <= #TCQ s_axis_tx_tdata;
          tvalid_prev  <= #TCQ s_axis_tx_tvalid;
          tkeep_prev   <= #TCQ s_axis_tx_tkeep;
          tlast_prev   <= #TCQ s_axis_tx_tlast;
          tuser_prev   <= #TCQ s_axis_tx_tuser;
        end
      end
    end

    // Create special buffer which locks in the proper value of TDATA depending
    // on whether the user is throttling or not. This buffer has three states:
    //
    //       HOLD state: TDATA maintains its current value
    //                   - the Block has throttled the PCIe block
    //   PREVIOUS state: the buffer provides the previous value on TDATA
    //                   - the Block has finished throttling, and is a little
    //                     behind the user
    //    CURRENT state: the buffer passes the current value on TDATA
    //                   - the Block is caught up and ready to receive the
    //                     latest data from the user
    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_tdata  <= #TCQ {C_DATA_WIDTH{1'b0}};
        reg_tvalid <= #TCQ 1'b0;
        reg_tkeep  <= #TCQ {KEEP_WIDTH{1'b0}};
        reg_tlast  <= #TCQ 1'b0;
        reg_tuser  <= #TCQ 4'h0;

        reg_tdst_rdy <= #TCQ 1'b0;
      end
      else begin
        reg_tdst_rdy <= #TCQ trn_tdst_rdy;

        if(!data_hold) begin
          // PREVIOUS state
          if(data_prev) begin
            reg_tdata  <= #TCQ tdata_prev;
            reg_tvalid <= #TCQ tvalid_prev;
            reg_tkeep  <= #TCQ tkeep_prev;
            reg_tlast  <= #TCQ tlast_prev;
            reg_tuser  <= #TCQ tuser_prev;
          end

          // CURRENT state
          else begin
            reg_tdata  <= #TCQ s_axis_tx_tdata;
            reg_tvalid <= #TCQ s_axis_tx_tvalid;
            reg_tkeep  <= #TCQ s_axis_tx_tkeep;
            reg_tlast  <= #TCQ s_axis_tx_tlast;
            reg_tuser  <= #TCQ s_axis_tx_tuser;
          end
        end
        // else HOLD state
      end
    end


    // Logic to instruct pipeline to hold its value
    assign data_hold = trn_tsrc_rdy && !trn_tdst_rdy;


    // Logic to instruct pipeline to use previous bus values. Always use
    // previous value after holding a value.
    always @(posedge user_clk) begin
      if(user_rst) begin
        data_prev <= #TCQ 1'b0;
      end
      else begin
        data_prev <= #TCQ data_hold;
      end
    end


    //------------------------------------------------------------------------//
    // Create trn_tsrc_rdy. If we're flushing the TRN hold trn_tsrc_rdy low.  //
    //------------------------------------------------------------------------//
    assign trn_tsrc_rdy = reg_tvalid && !disable_trn;


    //------------------------------------------------------------------------//
    // Create TREADY                                                          //
    //------------------------------------------------------------------------//
    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_tready <= #TCQ 1'b0;
      end
      else begin
        // If the link went down and we need to flush a packet in flight, hold
        // TREADY high
        if(flush_axi && !axi_end_packet) begin
          reg_tready <= #TCQ 1'b1;
        end

        // If the link is up, TREADY is as follows:
        //   TREADY = 1 when trn_tsrc_rdy == 0
        //      - While idle, keep the pipeline primed and ready for the next
        //        packet
        //
        //   TREADY = trn_tdst_rdy when trn_tsrc_rdy == 1
        //      - While in packet, throttle pipeline based on state of TRN
        else if(trn_lnk_up) begin
          reg_tready <= #TCQ trn_tdst_rdy || !trn_tsrc_rdy;
        end

        // If the link is down and we're not flushing a packet, hold TREADY low
        // wait for link to come back up
        else begin
          reg_tready <= #TCQ 1'b0;
        end
      end
    end

    assign s_axis_tx_tready = reg_tready;
  end


  //--------------------------------------------------------------------------//
  // Create flush_axi. This signal detects if the link goes down while the    //
  // AXI interface is in packet. In this situation, we need to flush the      //
  // packet through the AXI interface and discard it.                         //
  //--------------------------------------------------------------------------//
  always @(posedge user_clk) begin
    if(user_rst) begin
      flush_axi    <= #TCQ 1'b0;
    end
    else begin
      // If the AXI interface is in packet and the link goes down, purge it.
      if(axi_in_packet && !trn_lnk_up && !axi_end_packet) begin
        flush_axi <= #TCQ 1'b1;
      end

      // The packet is finished, so we're done flushing.
      else if(axi_end_packet) begin
        flush_axi <= #TCQ 1'b0;
      end
    end
  end
endgenerate

endmodule



`timescale 1ns/1ps
module model_ap2_tst_axi_basic_tx_thrtl_ctl #(
  parameter C_DATA_WIDTH = 128,           // RX/TX interface data width
  parameter C_FAMILY     = "X7",          // Targeted FPGA family
  parameter C_ROOT_PORT  = "FALSE",       // PCIe block is in root port mode
  parameter TCQ = 1                       // Clock to Q time
  ) (

  // AXI TX
  //-----------
  input  [C_DATA_WIDTH-1:0] s_axis_tx_tdata,         // TX data from user
  input                     s_axis_tx_tvalid,        // TX data is valid
  input               [3:0] s_axis_tx_tuser,         // TX user signals
  input                     s_axis_tx_tlast,         // TX data is last

  // User Misc.
  //-----------
  input                     user_turnoff_ok,         // Turnoff OK from user
  input                     user_tcfg_gnt,           // Send cfg OK from user

  // TRN TX
  //-----------
  input               [5:0] trn_tbuf_av,             // TX buffers available
  input                     trn_tdst_rdy,            // TX destination ready

  // TRN Misc.
  //-----------
  input                     trn_tcfg_req,            // TX config request
  output                    trn_tcfg_gnt,            // TX config grant
  input                     trn_lnk_up,              // PCIe link up

  // 7 Series/Virtex6 PM
  //-----------
  input               [2:0] cfg_pcie_link_state,     // Encoded PCIe link state

  // Virtex6 PM
  //-----------
  input                     cfg_pm_send_pme_to,      // PM send PME turnoff msg
  input               [1:0] cfg_pmcsr_powerstate,    // PMCSR power state
  input              [31:0] trn_rdllp_data,          // RX DLLP data
  input                     trn_rdllp_src_rdy,       // RX DLLP source ready

  // Virtex6/Spartan6 PM
  //-----------
  input                     cfg_to_turnoff,          // Turnoff request
  output reg                cfg_turnoff_ok,          // Turnoff grant

  // System
  //-----------
  output reg                tready_thrtl,            // TREADY to pipeline
  input                     user_clk,                // user clock from block
  input                     user_rst                 // user reset from block
);

// Thrtl user when TBUF hits this val
localparam TBUF_AV_MIN = (C_DATA_WIDTH == 128) ? 5 :
                                                   (C_DATA_WIDTH == 64) ? 1 : 0;

// Pause user when TBUF hits this val
localparam TBUF_AV_GAP = TBUF_AV_MIN + 1;

// GAP pause time - the latency from the time a packet is accepted on the TRN
// interface to the time trn_tbuf_av from the Block will decrement.
localparam TBUF_GAP_TIME = (C_DATA_WIDTH == 128) ? 4 : 1;

// Latency time from when tcfg_gnt is asserted to when PCIe block will throttle
localparam TCFG_LATENCY_TIME = 2'd2;

// Number of pipeline stages to delay trn_tcfg_gnt. For V6 128-bit only
localparam TCFG_GNT_PIPE_STAGES = 3;

// Throttle condition registers and constants
reg        lnk_up_thrtl;
wire       lnk_up_trig;
wire       lnk_up_exit;

reg        tbuf_av_min_thrtl;
wire       tbuf_av_min_trig;

reg        tbuf_av_gap_thrtl;
reg  [2:0] tbuf_gap_cnt;
wire       tbuf_av_gap_trig;
wire       tbuf_av_gap_exit;
wire       gap_trig_tlast;
wire       gap_trig_tcfg;
wire       gap_trig_decr;
reg  [5:0] tbuf_av_d;

reg        tcfg_req_thrtl;
reg  [1:0] tcfg_req_cnt;
reg        trn_tdst_rdy_d;
wire       tcfg_req_trig;
wire       tcfg_req_exit;
reg        tcfg_gnt_log;

wire       pre_throttle;
wire       reg_throttle;
wire       exit_crit;
reg        reg_tcfg_gnt;
reg        trn_tcfg_req_d;
reg        tcfg_gnt_pending;
wire       wire_to_turnoff;
reg        reg_turnoff_ok;

reg        tready_thrtl_mux;

localparam LINKSTATE_L0             = 3'b000;
localparam LINKSTATE_PPM_L1         = 3'b001;
localparam LINKSTATE_PPM_L1_TRANS   = 3'b101;
localparam LINKSTATE_PPM_L23R_TRANS = 3'b110;
localparam PM_ENTER_L1              = 8'h20;
localparam POWERSTATE_D0            = 2'b00;

reg        ppm_L1_thrtl;
wire       ppm_L1_trig;
wire       ppm_L1_exit;
reg  [2:0] cfg_pcie_link_state_d;
reg        trn_rdllp_src_rdy_d;

reg        ppm_L23_thrtl;
wire       ppm_L23_trig;
reg        cfg_turnoff_ok_pending;

reg        reg_tlast;

// Throttle control state machine states and registers
localparam IDLE       = 0;
localparam THROTTLE   = 1;
reg        cur_state;
reg        next_state;

reg        reg_axi_in_pkt;
wire       axi_in_pkt;
wire       axi_pkt_ending;
wire       axi_throttled;
wire       axi_thrtl_ok;
wire       tx_ecrc_pause;

//----------------------------------------------------------------------------//
// THROTTLE REASON: PCIe link is down                                         //
//   - When to throttle: trn_lnk_up deasserted                                //
//   - When to stop: trn_tdst_rdy assesrted                                   //
//----------------------------------------------------------------------------//
assign lnk_up_trig = !trn_lnk_up;
assign lnk_up_exit = trn_tdst_rdy;

always @(posedge user_clk) begin
  if(user_rst) begin
    lnk_up_thrtl <= #TCQ 1'b1;
  end
  else begin
    if(lnk_up_trig) begin
      lnk_up_thrtl <= #TCQ 1'b1;
    end
    else if(lnk_up_exit) begin
      lnk_up_thrtl <= #TCQ 1'b0;
    end
  end
end


//----------------------------------------------------------------------------//
// THROTTLE REASON: Transmit buffers depleted                                 //
//   - When to throttle: trn_tbuf_av falls to 0                               //
//   - When to stop: trn_tbuf_av rises above 0 again                          //
//----------------------------------------------------------------------------//
assign tbuf_av_min_trig = (trn_tbuf_av <= TBUF_AV_MIN);

always @(posedge user_clk) begin
  if(user_rst) begin
    tbuf_av_min_thrtl <= #TCQ 1'b0;
  end
  else begin
    if(tbuf_av_min_trig) begin
      tbuf_av_min_thrtl <= #TCQ 1'b1;
    end

    // The exit condition for tbuf_av_min_thrtl is !tbuf_av_min_trig
    else begin
      tbuf_av_min_thrtl <= #TCQ 1'b0;
    end
  end
end


//----------------------------------------------------------------------------//
// THROTTLE REASON: Transmit buffers getting low                              //
//   - When to throttle: trn_tbuf_av falls below "gap" threshold TBUF_AV_GAP  //
//   - When to stop: after TBUF_GAP_TIME cycles elapse                        //
//                                                                            //
// If we're about to run out of transmit buffers, throttle the user for a     //
// few clock cycles to give the PCIe block time to catch up. This is          //
// needed to compensate for latency in decrementing trn_tbuf_av in the PCIe   //
// Block transmit path.                                                       //
//----------------------------------------------------------------------------//

// Detect two different scenarios for buffers getting low:
// 1) If we see a TLAST. a new packet has been inserted into the buffer, and
//    we need to pause and let that packet "soak in"
assign gap_trig_tlast = (trn_tbuf_av <= TBUF_AV_GAP) &&
                            s_axis_tx_tvalid && tready_thrtl && s_axis_tx_tlast;

// 2) Any time tbug_avail decrements to the TBUF_AV_GAP threshold, we need to
//    pause and make sure no other packets are about to soak in and cause the
//    buffer availability to drop further.
assign gap_trig_decr  = (trn_tbuf_av == (TBUF_AV_GAP)) &&
                                                 (tbuf_av_d == (TBUF_AV_GAP+1));

assign gap_trig_tcfg  = (tcfg_req_thrtl && tcfg_req_exit);
assign tbuf_av_gap_trig = gap_trig_tlast || gap_trig_decr || gap_trig_tcfg;
assign tbuf_av_gap_exit = (tbuf_gap_cnt == 0);

always @(posedge user_clk) begin
  if(user_rst) begin
    tbuf_av_gap_thrtl <= #TCQ 1'b0;
    tbuf_gap_cnt      <= #TCQ 3'h0;
    tbuf_av_d         <= #TCQ 6'h00;
  end
  else begin
    if(tbuf_av_gap_trig) begin
      tbuf_av_gap_thrtl <= #TCQ 1'b1;
    end
    else if(tbuf_av_gap_exit) begin
      tbuf_av_gap_thrtl <= #TCQ 1'b0;
    end

    // tbuf gap counter:
    // This logic controls the length of the throttle condition when tbufs are
    // getting low.
    if(tbuf_av_gap_thrtl && (cur_state == THROTTLE)) begin
      if(tbuf_gap_cnt > 0) begin
        tbuf_gap_cnt <= #TCQ tbuf_gap_cnt - 3'd1;
      end
    end
    else begin
      tbuf_gap_cnt <= #TCQ TBUF_GAP_TIME;
    end

    tbuf_av_d <= #TCQ trn_tbuf_av;
  end
end


//----------------------------------------------------------------------------//
// THROTTLE REASON: Block needs to send a CFG response                        //
//   - When to throttle: trn_tcfg_req and user_tcfg_gnt asserted              //
//   - When to stop: after trn_tdst_rdy transitions to unasserted             //
//                                                                            //
// If the block needs to send a response to a CFG packet, this will cause     //
// the subsequent deassertion of trn_tdst_rdy. When the user design permits,  //
// grant permission to the block to service request and throttle the user.    //
//----------------------------------------------------------------------------//
assign tcfg_req_trig = trn_tcfg_req && reg_tcfg_gnt;
assign tcfg_req_exit = (tcfg_req_cnt == 2'd0) && !trn_tdst_rdy_d &&
                                                                   trn_tdst_rdy;
always @(posedge user_clk) begin
  if(user_rst) begin
    tcfg_req_thrtl   <= #TCQ 1'b0;
    trn_tcfg_req_d   <= #TCQ 1'b0;
    trn_tdst_rdy_d   <= #TCQ 1'b1;
    reg_tcfg_gnt     <= #TCQ 1'b0;
    tcfg_req_cnt     <= #TCQ 2'd0;
    tcfg_gnt_pending <= #TCQ 1'b0;
  end
  else begin
    if(tcfg_req_trig) begin
      tcfg_req_thrtl <= #TCQ 1'b1;
    end
    else if(tcfg_req_exit) begin
      tcfg_req_thrtl <= #TCQ 1'b0;
    end

    // We need to wait the appropriate amount of time for the tcfg_gnt to
    // "sink in" to the PCIe block. After that, we know that the PCIe block will
    // not reassert trn_tdst_rdy until the CFG request has been serviced. If a
    // new request is being service (tcfg_gnt_log == 1), then reset the timer.
    if((trn_tcfg_req && !trn_tcfg_req_d) || tcfg_gnt_pending) begin
      tcfg_req_cnt <= #TCQ TCFG_LATENCY_TIME;
    end
    else begin
      if(tcfg_req_cnt > 0) begin
        tcfg_req_cnt <= #TCQ tcfg_req_cnt - 2'd1;
      end
    end

    // Make sure tcfg_gnt_log pulses once for one clock cycle for every
    // cfg packet request.
    if(trn_tcfg_req && !trn_tcfg_req_d) begin
      tcfg_gnt_pending <= #TCQ 1'b1;
    end
    else if(tcfg_gnt_log) begin
      tcfg_gnt_pending <= #TCQ 1'b0;
    end

    trn_tcfg_req_d <= #TCQ trn_tcfg_req;
    trn_tdst_rdy_d <= #TCQ trn_tdst_rdy;
    reg_tcfg_gnt   <= #TCQ user_tcfg_gnt;
  end
end


//----------------------------------------------------------------------------//
// THROTTLE REASON: Block needs to transition to low power state PPM L1       //
//   - When to throttle: appropriate low power state signal asserted          //
//     (architecture dependent)                                               //
//   - When to stop: cfg_pcie_link_state goes to proper value (C_ROOT_PORT    //
//     dependent)                                                             //
//                                                                            //
// If the block needs to transition to PM state PPM L1, we need to finish     //
// up what we're doing and throttle immediately.                              //
//----------------------------------------------------------------------------//
generate
  // PPM L1 signals for 7 Series in RC mode
  if((C_FAMILY == "X7") && (C_ROOT_PORT == "TRUE")) begin : x7_L1_thrtl_rp
    assign ppm_L1_trig = (cfg_pcie_link_state_d == LINKSTATE_L0) &&
                           (cfg_pcie_link_state == LINKSTATE_PPM_L1_TRANS);
    assign ppm_L1_exit = cfg_pcie_link_state == LINKSTATE_PPM_L1;
  end

  // PPM L1 signals for 7 Series in EP mode
  else if((C_FAMILY == "X7") && (C_ROOT_PORT == "FALSE")) begin : x7_L1_thrtl_ep
    assign ppm_L1_trig = (cfg_pcie_link_state_d == LINKSTATE_L0) &&
                           (cfg_pcie_link_state == LINKSTATE_PPM_L1_TRANS);
    assign ppm_L1_exit = cfg_pcie_link_state == LINKSTATE_L0;
  end

  // PPM L1 signals for V6 in RC mode
  else if((C_FAMILY == "V6") && (C_ROOT_PORT == "TRUE")) begin : v6_L1_thrtl_rp
    assign ppm_L1_trig = (trn_rdllp_data[31:24] == PM_ENTER_L1) &&
                                      trn_rdllp_src_rdy && !trn_rdllp_src_rdy_d;
    assign ppm_L1_exit = cfg_pcie_link_state == LINKSTATE_PPM_L1;
  end

  // PPM L1 signals for V6 in EP mode
  else if((C_FAMILY == "V6") && (C_ROOT_PORT == "FALSE")) begin : v6_L1_thrtl_ep
    assign ppm_L1_trig = (cfg_pmcsr_powerstate != POWERSTATE_D0);
    assign ppm_L1_exit = cfg_pcie_link_state == LINKSTATE_L0;
  end

  // PPM L1 detection not supported for S6
  else begin : s6_L1_thrtl
    assign ppm_L1_trig = 1'b0;
    assign ppm_L1_exit = 1'b1;
  end
endgenerate

always @(posedge user_clk) begin
  if(user_rst) begin
    ppm_L1_thrtl          <= #TCQ 1'b0;
    cfg_pcie_link_state_d <= #TCQ 3'b0;
    trn_rdllp_src_rdy_d   <= #TCQ 1'b0;
  end
  else begin
    if(ppm_L1_trig) begin
      ppm_L1_thrtl <= #TCQ 1'b1;
    end
    else if(ppm_L1_exit) begin
      ppm_L1_thrtl <= #TCQ 1'b0;
    end
    cfg_pcie_link_state_d <= #TCQ cfg_pcie_link_state;
    trn_rdllp_src_rdy_d   <= #TCQ trn_rdllp_src_rdy;
  end
end


//----------------------------------------------------------------------------//
// THROTTLE REASON: Block needs to transition to low power state PPM L2/3     //
//   - When to throttle: appropriate PM signal indicates a transition to      //
//     L2/3 is pending or in progress (family and role dependent)             //
//   - When to stop: never (the only path out of L2/3 is a full reset)        //
//                                                                            //
// If the block needs to transition to PM state PPM L2/3, we need to finish   //
// up what we're doing and throttle when the user gives permission.           //
//----------------------------------------------------------------------------//
generate
  // PPM L2/3 signals for 7 Series in RC mode
  if((C_FAMILY == "X7") && (C_ROOT_PORT == "TRUE")) begin : x7_L23_thrtl_rp
    assign ppm_L23_trig = (cfg_pcie_link_state_d == LINKSTATE_PPM_L23R_TRANS);
    assign wire_to_turnoff = 1'b0;
  end

  // PPM L2/3 signals for V6 in RC mode
  else if((C_FAMILY == "V6") && (C_ROOT_PORT == "TRUE")) begin : v6_L23_thrtl_rp
    assign ppm_L23_trig = cfg_pm_send_pme_to;
    assign wire_to_turnoff = 1'b0;
  end

  // PPM L2/3 signals in EP mode
  else begin : L23_thrtl_ep
    assign ppm_L23_trig = wire_to_turnoff && reg_turnoff_ok;

    // PPM L2/3 signals for 7 Series in EP mode
    // For 7 Series, cfg_to_turnoff pulses once when a turnoff request is
    // outstanding, so we need a "sticky" register that grabs the request.
    if(C_FAMILY == "X7") begin : x7_L23_thrtl_ep
      reg reg_to_turnoff;

      always @(posedge user_clk) begin
        if(user_rst) begin
          reg_to_turnoff <= #TCQ 1'b0;
        end
        else begin
          if(cfg_to_turnoff) begin
            reg_to_turnoff <= #TCQ 1'b1;
          end
        end
      end

      assign wire_to_turnoff = reg_to_turnoff;
    end

    // PPM L2/3 signals for V6/S6 in EP mode
    // In V6 and S6, the to_turnoff signal asserts and remains asserted until
    // turnoff_ok is asserted, so a sticky reg is not necessary.
    else begin : v6_s6_L23_thrtl_ep
      assign wire_to_turnoff = cfg_to_turnoff;
    end

    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_turnoff_ok <= #TCQ 1'b0;
      end
      else begin
        reg_turnoff_ok <= #TCQ user_turnoff_ok;
      end
    end
  end
endgenerate

always @(posedge user_clk) begin
  if(user_rst) begin
    ppm_L23_thrtl   <= #TCQ 1'b0;
    cfg_turnoff_ok_pending <= #TCQ 1'b0;
  end
  else begin
    if(ppm_L23_trig) begin
      ppm_L23_thrtl <= #TCQ 1'b1;
    end

    // Make sure cfg_turnoff_ok pulses once for one clock cycle for every
    // turnoff request.
    if(ppm_L23_trig && !ppm_L23_thrtl) begin
      cfg_turnoff_ok_pending <= #TCQ 1'b1;
    end
    else if(cfg_turnoff_ok) begin
      cfg_turnoff_ok_pending <= #TCQ 1'b0;
    end
  end
end


//----------------------------------------------------------------------------//
// Create axi_thrtl_ok. This signal determines if it's OK to throttle the     //
// user design on the AXI interface. Since TREADY is registered, this signal  //
// needs to assert on the cycle ~before~ we actually intend to throttle.      //
// The only time it's OK to throttle when TVALID is asserted is on the first  //
// beat of a new packet. Therefore, assert axi_thrtl_ok if one of the         //
// is true:                                                                   //
//    1) The user is not in a packet and is not starting one                  //
//    2) The user is just finishing a packet                                  //
//    3) We're already throttled, so it's OK to continue throttling           //
//----------------------------------------------------------------------------//
always @(posedge user_clk) begin
  if(user_rst) begin
    reg_axi_in_pkt <= #TCQ 1'b0;
  end
  else begin
    if(s_axis_tx_tvalid && s_axis_tx_tlast) begin
      reg_axi_in_pkt <= #TCQ 1'b0;
    end
    else if(tready_thrtl && s_axis_tx_tvalid) begin
      reg_axi_in_pkt <= #TCQ 1'b1;
    end
  end
end

assign axi_in_pkt     = s_axis_tx_tvalid || reg_axi_in_pkt;
assign axi_pkt_ending = s_axis_tx_tvalid && s_axis_tx_tlast;
assign axi_throttled  = !tready_thrtl;
assign axi_thrtl_ok   = !axi_in_pkt || axi_pkt_ending || axi_throttled;


//----------------------------------------------------------------------------//
// Throttle CTL State Machine:                                                //
// Throttle user design when a throttle trigger (or triggers) occur.          //
// Keep user throttled until all exit criteria have been met.                 //
//----------------------------------------------------------------------------//

// Immediate throttle signal. Used to "pounce" on a throttle opportunity when
// we're seeking one
assign pre_throttle = tbuf_av_min_trig || tbuf_av_gap_trig || lnk_up_trig
                                || tcfg_req_trig || ppm_L1_trig || ppm_L23_trig;


// Registered throttle signals. Used to control throttle state machine
assign reg_throttle = tbuf_av_min_thrtl || tbuf_av_gap_thrtl || lnk_up_thrtl
                             || tcfg_req_thrtl || ppm_L1_thrtl || ppm_L23_thrtl;

assign exit_crit = !tbuf_av_min_thrtl && !tbuf_av_gap_thrtl && !lnk_up_thrtl
                          && !tcfg_req_thrtl && !ppm_L1_thrtl && !ppm_L23_thrtl;

always @(*) begin
  case(cur_state)
    // IDLE: in this state we're waiting for a trigger event to occur. As
    // soon as an event occurs and the user isn't transmitting a packet, we
    // throttle the PCIe block and the user and next state is THROTTLE.
    IDLE: begin
      if(reg_throttle && axi_thrtl_ok) begin
        // Throttle user
        tready_thrtl_mux = 1'b0;
        next_state       = THROTTLE;

        // Assert appropriate grant signal depending on the throttle type.
        if(tcfg_req_thrtl) begin
          tcfg_gnt_log   = 1'b1;   // For cfg request, grant the request
          cfg_turnoff_ok = 1'b0;   //
        end
        else if(ppm_L23_thrtl) begin
          tcfg_gnt_log   = 1'b0;   //
          cfg_turnoff_ok = 1'b1;   // For PM request, permit transition
        end
        else begin
          tcfg_gnt_log   = 1'b0;   // Otherwise do nothing
          cfg_turnoff_ok = 1'b0;   //
        end
      end

      // If there's not throttle event, do nothing
      else begin
        // Throttle user as soon as possible
        tready_thrtl_mux = !(axi_thrtl_ok && pre_throttle);
        next_state       = IDLE;

        tcfg_gnt_log     = 1'b0;
        cfg_turnoff_ok   = 1'b0;
      end
    end

    // THROTTLE: in this state the user is throttle and we're waiting for
    // exit criteria, which tells us that the throttle event is over. When
    // the exit criteria is satisfied, de-throttle the user and next state
    // is IDLE.
    THROTTLE: begin
      if(exit_crit) begin
        // Dethrottle user
        tready_thrtl_mux = !pre_throttle;
        next_state       = IDLE;
      end
      else begin
        // Throttle user
        tready_thrtl_mux = 1'b0;
        next_state       = THROTTLE;
      end

      // Assert appropriate grant signal depending on the throttle type.
      if(tcfg_req_thrtl && tcfg_gnt_pending) begin
        tcfg_gnt_log   = 1'b1;   // For cfg request, grant the request
        cfg_turnoff_ok = 1'b0;   //
      end
      else if(cfg_turnoff_ok_pending) begin
        tcfg_gnt_log   = 1'b0;   //
        cfg_turnoff_ok = 1'b1;   // For PM request, permit transition
      end
      else begin
        tcfg_gnt_log   = 1'b0;   // Otherwise do nothing
        cfg_turnoff_ok = 1'b0;   //
      end
    end

    default: begin
      tready_thrtl_mux = 1'b0;
      next_state       = IDLE;
      tcfg_gnt_log     = 1'b0;
      cfg_turnoff_ok   = 1'b0;
    end
  endcase
end

// Synchronous logic
always @(posedge user_clk) begin
  if(user_rst) begin
    // Throttle user by default until link comes up
    cur_state        <= #TCQ THROTTLE;

    reg_tlast        <= #TCQ 1'b0;

    tready_thrtl     <= #TCQ 1'b0;
  end
  else begin
    cur_state        <= #TCQ next_state;

    tready_thrtl     <= #TCQ tready_thrtl_mux && !tx_ecrc_pause;
    reg_tlast        <= #TCQ s_axis_tx_tlast;
  end
end

// For X7, the PCIe block will generate the ECRC for a packet if trn_tecrc_gen
// is asserted at SOF. In this case, the Block needs an extra data beat to
// calculate the ECRC, but only if the following conditions are met:
//  1) there is no empty DWORDS at the end of the packet
//     (i.e. packet length % C_DATA_WIDTH == 0)
//
//  2) There isn't a ECRC in the TLP already, as indicated by the TD bit in the
//     TLP header
//
// If both conditions are met, the Block will stall the TRN interface for one
// data beat after EOF. We need to predict this stall and preemptively stall the
// User for one beat.
generate
  if(C_FAMILY == "X7") begin : ecrc_pause_enabled
    wire        tx_ecrc_pkt;
    reg         reg_tx_ecrc_pkt;

    wire  [1:0] packet_fmt;
    wire        packet_td;
    wire  [2:0] header_len;
    wire  [9:0] payload_len;
    wire [13:0] packet_len;
    wire        pause_needed;

    // Grab necessary packet fields
    assign packet_fmt  = s_axis_tx_tdata[30:29];
    assign packet_td   = s_axis_tx_tdata[15];

    // Calculate total packet length
    assign header_len  = packet_fmt[0] ? 3'd4 : 3'd3;
    assign payload_len = packet_fmt[1] ? s_axis_tx_tdata[9:0] : 10'h0;
    assign packet_len  = {10'h000, header_len} + {4'h0, payload_len};


    // Determine if packet a ECRC pause is needed
    if(C_DATA_WIDTH == 128) begin : packet_len_check_128
      assign pause_needed = (packet_len[1:0] == 2'b00) && !packet_td;
    end
    else begin : packet_len_check_64
      assign pause_needed = (packet_len[0] == 1'b0) && !packet_td;
    end


    // Create flag to alert TX pipeline to insert a stall
    assign tx_ecrc_pkt = s_axis_tx_tuser[0] && pause_needed &&
                            tready_thrtl && s_axis_tx_tvalid && !reg_axi_in_pkt;

    always @(posedge user_clk) begin
      if(user_rst) begin
        reg_tx_ecrc_pkt <= #TCQ 1'b0;
      end
      else begin
        if(tx_ecrc_pkt && !s_axis_tx_tlast) begin
          reg_tx_ecrc_pkt <= #TCQ 1'b1;
        end
        else if(tready_thrtl && s_axis_tx_tvalid && s_axis_tx_tlast) begin
          reg_tx_ecrc_pkt <= #TCQ 1'b0;
        end
      end
    end


    // Insert the stall now
    assign tx_ecrc_pause = ((tx_ecrc_pkt || reg_tx_ecrc_pkt) &&
                           s_axis_tx_tlast && s_axis_tx_tvalid && tready_thrtl);

  end
  else begin : ecrc_pause_disabled
    assign tx_ecrc_pause = 1'b0;
  end
endgenerate


// Logic for 128-bit single cycle bug fix.
// This tcfg_gnt pipeline addresses an issue with 128-bit V6 designs where a
// single cycle packet transmitted simultaneously with an assertion of tcfg_gnt
// from AXI Basic causes the packet to be dropped. The packet drop occurs
// because the 128-bit shim doesn't know about the tcfg_req/gnt, and therefor
// isn't expecting trn_tdst_rdy to go low. Since the 128-bit shim does throttle
// prediction just as we do, it ignores the value of trn_tdst_rdy, and
// ultimately drops the packet when transmitting the packet to the block.
generate
  if(C_DATA_WIDTH == 128 && C_FAMILY == "V6") begin : tcfg_gnt_pipeline
    genvar stage;
    reg tcfg_gnt_pipe [TCFG_GNT_PIPE_STAGES:0];

    // Create a configurable depth FF delay pipeline
    for(stage = 0; stage < TCFG_GNT_PIPE_STAGES; stage = stage + 1)
    begin : tcfg_gnt_pipeline_stage

      always @(posedge user_clk) begin
        if(user_rst) begin
          tcfg_gnt_pipe[stage] <= #TCQ 1'b0;
        end
        else begin
          // For stage 0, insert the actual tcfg_gnt signal from logic
          if(stage == 0) begin
            tcfg_gnt_pipe[stage] <= #TCQ tcfg_gnt_log;
          end

          // For stages 1+, chain together
          else begin
            tcfg_gnt_pipe[stage] <= #TCQ tcfg_gnt_pipe[stage - 1];
          end
        end
      end

      // tcfg_gnt output to block assigned the last pipeline stage
      assign trn_tcfg_gnt = tcfg_gnt_pipe[TCFG_GNT_PIPE_STAGES-1];
    end
  end
  else begin : tcfg_gnt_no_pipeline

    // For all other architectures, no pipeline delay needed for tcfg_gnt
    assign trn_tcfg_gnt = tcfg_gnt_log;
  end
endgenerate

endmodule


`timescale 1ns/1ps
module model_ap2_tst_pcie_7x # (
  // PCIE_2_1 params
  parameter [11:0] AER_BASE_PTR = 12'h140,
  parameter        AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter        AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [15:0] AER_CAP_ID = 16'h0001,
  parameter        AER_CAP_MULTIHEADER = "FALSE",
  parameter [11:0] AER_CAP_NEXTPTR = 12'h178,
  parameter        AER_CAP_ON = "FALSE",
  parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000,
  parameter        AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE",
  parameter [3:0]  AER_CAP_VERSION = 4'h1,
  parameter        ALLOW_X8_GEN2 = "FALSE",
  parameter [31:0] BAR0 = 32'hFFFFFF00,
  parameter [31:0] BAR1 = 32'hFFFF0000,
  parameter [31:0] BAR2 = 32'hFFFF000C,
  parameter [31:0] BAR3 = 32'hFFFFFFFF,
  parameter [31:0] BAR4 = 32'h00000000,
  parameter [31:0] BAR5 = 32'h00000000,
  parameter [7:0]  CAPABILITIES_PTR = 8'h40,
  parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000,
  parameter        CFG_ECRC_ERR_CPLSTAT = 0,
  parameter [23:0] CLASS_CODE = 24'h000000,
  parameter        CMD_INTX_IMPLEMENTED = "TRUE",
  parameter        CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE",
  parameter [3:0]  CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0,
  parameter [6:0]  CRM_MODULE_RSTS = 7'h00,
  parameter        C_DATA_WIDTH = 64,
  parameter        REM_WIDTH = (C_DATA_WIDTH == 128) ? 2 : 1,
  parameter        KEEP_WIDTH = C_DATA_WIDTH / 8,
  parameter        DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE",
  parameter        DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE",
  parameter [1:0]  DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0,
  parameter        DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE",
  parameter [1:0]  DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0,
  parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE",
  parameter        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE",
  parameter        integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0,
  parameter        integer DEV_CAP_ENDPOINT_L1_LATENCY = 0,
  parameter        DEV_CAP_EXT_TAG_SUPPORTED = "TRUE",
  parameter        DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE",
  parameter        integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2,
  parameter        integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0,
  parameter        DEV_CAP_ROLE_BASED_ERROR = "TRUE",
  parameter        integer DEV_CAP_RSVD_14_12 = 0,
  parameter        integer DEV_CAP_RSVD_17_16 = 0,
  parameter        integer DEV_CAP_RSVD_31_29 = 0,
  parameter        DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE",
  parameter        DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE",
  parameter        DISABLE_ASPM_L1_TIMER = "FALSE",
  parameter        DISABLE_BAR_FILTERING = "FALSE",
  parameter        DISABLE_ERR_MSG = "FALSE",
  parameter        DISABLE_ID_CHECK = "FALSE",
  parameter        DISABLE_LANE_REVERSAL = "FALSE",
  parameter        DISABLE_LOCKED_FILTER = "FALSE",
  parameter        DISABLE_PPM_FILTER = "FALSE",
  parameter        DISABLE_RX_POISONED_RESP = "FALSE",
  parameter        DISABLE_RX_TC_FILTER = "FALSE",
  parameter        DISABLE_SCRAMBLING = "FALSE",
  parameter [7:0]  DNSTREAM_LINK_NUM = 8'h00,
  parameter [11:0] DSN_BASE_PTR = 12'h100,
  parameter [15:0] DSN_CAP_ID = 16'h0003,
  parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C,
  parameter        DSN_CAP_ON = "TRUE",
  parameter [3:0]  DSN_CAP_VERSION = 4'h1,
  parameter [10:0] ENABLE_MSG_ROUTE = 11'h000,
  parameter        ENABLE_RX_TD_ECRC_TRIM = "FALSE",
  parameter        ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE",
  parameter        ENTER_RVRY_EI_L0 = "TRUE",
  parameter        EXIT_LOOPBACK_ON_EI = "TRUE",
  parameter [31:0] EXPANSION_ROM = 32'hFFFFF001,
  parameter [5:0]  EXT_CFG_CAP_PTR = 6'h3F,
  parameter [9:0]  EXT_CFG_XP_CAP_PTR = 10'h3FF,
  parameter [7:0]  HEADER_TYPE = 8'h00,
  parameter [4:0]  INFER_EI = 5'h00,
  parameter [7:0]  INTERRUPT_PIN = 8'h01,
  parameter        INTERRUPT_STAT_AUTO = "TRUE",
  parameter        IS_SWITCH = "FALSE",
  parameter [9:0]  LAST_CONFIG_DWORD = 10'h3FF,
  parameter        LINK_CAP_ASPM_OPTIONALITY = "TRUE",
  parameter        integer LINK_CAP_ASPM_SUPPORT = 1,
  parameter        LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE",
  parameter        LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE",
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7,
  parameter        integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7,
  parameter        integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7,
  parameter        LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE",
  parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,
  parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,
  parameter        integer LINK_CAP_RSVD_23 = 0,
  parameter        LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE",
  parameter        integer LINK_CONTROL_RCB = 0,
  parameter        LINK_CTRL2_DEEMPHASIS = "FALSE",
  parameter        LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE",
  parameter [3:0]  LINK_CTRL2_TARGET_LINK_SPEED = 4'h2,
  parameter        LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE",
  parameter [14:0] LL_ACK_TIMEOUT = 15'h0000,
  parameter        LL_ACK_TIMEOUT_EN = "FALSE",
  parameter        integer LL_ACK_TIMEOUT_FUNC = 0,
  parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000,
  parameter        LL_REPLAY_TIMEOUT_EN = "FALSE",
  parameter        integer LL_REPLAY_TIMEOUT_FUNC = 0,
  parameter [5:0]  LTSSM_MAX_LINK_WIDTH = 6'h01,
  parameter        MPS_FORCE = "FALSE",
  parameter [7:0]  MSIX_BASE_PTR = 8'h9C,
  parameter [7:0]  MSIX_CAP_ID = 8'h11,
  parameter [7:0]  MSIX_CAP_NEXTPTR = 8'h00,
  parameter        MSIX_CAP_ON = "FALSE",
  parameter        integer MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter        integer MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter [7:0]  MSI_BASE_PTR = 8'h48,
  parameter        MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE",
  parameter [7:0]  MSI_CAP_ID = 8'h05,
  parameter        integer MSI_CAP_MULTIMSGCAP = 0,
  parameter        integer MSI_CAP_MULTIMSG_EXTENSION = 0,
  parameter [7:0]  MSI_CAP_NEXTPTR = 8'h60,
  parameter        MSI_CAP_ON = "FALSE",
  parameter        MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE",
  parameter        integer N_FTS_COMCLK_GEN1 = 255,
  parameter        integer N_FTS_COMCLK_GEN2 = 255,
  parameter        integer N_FTS_GEN1 = 255,
  parameter        integer N_FTS_GEN2 = 255,
  parameter [7:0]  PCIE_BASE_PTR = 8'h60,
  parameter [7:0]  PCIE_CAP_CAPABILITY_ID = 8'h10,
  parameter [3:0]  PCIE_CAP_CAPABILITY_VERSION = 4'h2,
  parameter [3:0]  PCIE_CAP_DEVICE_PORT_TYPE = 4'h0,
  parameter [7:0]  PCIE_CAP_NEXTPTR = 8'h9C,
  parameter        PCIE_CAP_ON = "TRUE",
  parameter        integer PCIE_CAP_RSVD_15_14 = 0,
  parameter        PCIE_CAP_SLOT_IMPLEMENTED = "FALSE",
  parameter        integer PCIE_REVISION = 2,
  parameter        integer PL_AUTO_CONFIG = 0,
  parameter        PL_FAST_TRAIN = "FALSE",
  parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000,
  parameter        PM_ASPML0S_TIMEOUT_EN = "FALSE",
  parameter        integer PM_ASPML0S_TIMEOUT_FUNC = 0,
  parameter        PM_ASPM_FASTEXIT = "FALSE",
  parameter [7:0]  PM_BASE_PTR = 8'h40,
  parameter        integer PM_CAP_AUXCURRENT = 0,
  parameter        PM_CAP_D1SUPPORT = "TRUE",
  parameter        PM_CAP_D2SUPPORT = "TRUE",
  parameter        PM_CAP_DSI = "FALSE",
  parameter [7:0]  PM_CAP_ID = 8'h01,
  parameter [7:0]  PM_CAP_NEXTPTR = 8'h48,
  parameter        PM_CAP_ON = "TRUE",
  parameter [4:0]  PM_CAP_PMESUPPORT = 5'h0F,
  parameter        PM_CAP_PME_CLOCK = "FALSE",
  parameter        integer PM_CAP_RSVD_04 = 0,
  parameter        integer PM_CAP_VERSION = 3,
  parameter        PM_CSR_B2B3 = "FALSE",
  parameter        PM_CSR_BPCCEN = "FALSE",
  parameter        PM_CSR_NOSOFTRST = "TRUE",
  parameter [7:0]  PM_DATA0 = 8'h01,
  parameter [7:0]  PM_DATA1 = 8'h01,
  parameter [7:0]  PM_DATA2 = 8'h01,
  parameter [7:0]  PM_DATA3 = 8'h01,
  parameter [7:0]  PM_DATA4 = 8'h01,
  parameter [7:0]  PM_DATA5 = 8'h01,
  parameter [7:0]  PM_DATA6 = 8'h01,
  parameter [7:0]  PM_DATA7 = 8'h01,
  parameter [1:0]  PM_DATA_SCALE0 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE1 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE2 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE3 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE4 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE5 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE6 = 2'h1,
  parameter [1:0]  PM_DATA_SCALE7 = 2'h1,
  parameter        PM_MF = "FALSE",
  parameter [11:0] RBAR_BASE_PTR = 12'h178,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00,
  parameter [4:0]  RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00,
  parameter [15:0] RBAR_CAP_ID = 16'h0015,
  parameter [2:0]  RBAR_CAP_INDEX0 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX1 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX2 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX3 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX4 = 3'h0,
  parameter [2:0]  RBAR_CAP_INDEX5 = 3'h0,
  parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000,
  parameter        RBAR_CAP_ON = "FALSE",
  parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000,
  parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000,
  parameter [3:0]  RBAR_CAP_VERSION = 4'h1,
  parameter [2:0]  RBAR_NUM = 3'h1,
  parameter        integer RECRC_CHK = 0,
  parameter        RECRC_CHK_TRIM = "FALSE",
  parameter        ROOT_CAP_CRS_SW_VISIBILITY = "FALSE",
  parameter [1:0]  RP_AUTO_SPD = 2'h1,
  parameter [4:0]  RP_AUTO_SPD_LOOPCNT = 5'h1f,
  parameter        SELECT_DLL_IF = "FALSE",
  parameter        SIM_VERSION = "1.0",
  parameter        SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE",
  parameter        SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE",
  parameter        SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE",
  parameter        SLOT_CAP_HOTPLUG_CAPABLE = "FALSE",
  parameter        SLOT_CAP_HOTPLUG_SURPRISE = "FALSE",
  parameter        SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE",
  parameter        SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE",
  parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000,
  parameter        SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE",
  parameter        SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE",
  parameter        integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0,
  parameter [7:0]  SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00,
  parameter        integer SPARE_BIT0 = 0,
  parameter        integer SPARE_BIT1 = 0,
  parameter        integer SPARE_BIT2 = 0,
  parameter        integer SPARE_BIT3 = 0,
  parameter        integer SPARE_BIT4 = 0,
  parameter        integer SPARE_BIT5 = 0,
  parameter        integer SPARE_BIT6 = 0,
  parameter        integer SPARE_BIT7 = 0,
  parameter        integer SPARE_BIT8 = 0,
  parameter [7:0]  SPARE_BYTE0 = 8'h00,
  parameter [7:0]  SPARE_BYTE1 = 8'h00,
  parameter [7:0]  SPARE_BYTE2 = 8'h00,
  parameter [7:0]  SPARE_BYTE3 = 8'h00,
  parameter [31:0] SPARE_WORD0 = 32'h00000000,
  parameter [31:0] SPARE_WORD1 = 32'h00000000,
  parameter [31:0] SPARE_WORD2 = 32'h00000000,
  parameter [31:0] SPARE_WORD3 = 32'h00000000,
  parameter        SSL_MESSAGE_AUTO = "FALSE",
  parameter        TECRC_EP_INV = "FALSE",
  parameter        TL_RBYPASS = "FALSE",
  parameter        integer TL_RX_RAM_RADDR_LATENCY = 0,
  parameter        integer TL_RX_RAM_RDATA_LATENCY = 2,
  parameter        integer TL_RX_RAM_WRITE_LATENCY = 0,
  parameter        TL_TFC_DISABLE = "FALSE",
  parameter        TL_TX_CHECKS_DISABLE = "FALSE",
  parameter        integer TL_TX_RAM_RADDR_LATENCY = 0,
  parameter        integer TL_TX_RAM_RDATA_LATENCY = 2,
  parameter        integer TL_TX_RAM_WRITE_LATENCY = 0,
  parameter        TRN_DW = "FALSE",
  parameter        TRN_NP_FC = "FALSE",
  parameter        UPCONFIG_CAPABLE = "TRUE",
  parameter        UPSTREAM_FACING = "TRUE",
  parameter        UR_ATOMIC = "TRUE",
  parameter        UR_CFG1 = "TRUE",
  parameter        UR_INV_REQ = "TRUE",
  parameter        UR_PRS_RESPONSE = "TRUE",
  parameter        USER_CLK2_DIV2 = "FALSE",
  parameter        integer USER_CLK_FREQ = 3,
  parameter        USE_RID_PINS = "FALSE",
  parameter        VC0_CPL_INFINITE = "TRUE",
  parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF,
  parameter        integer VC0_TOTAL_CREDITS_CD = 127,
  parameter        integer VC0_TOTAL_CREDITS_CH = 31,
  parameter        integer VC0_TOTAL_CREDITS_NPD = 24,
  parameter        integer VC0_TOTAL_CREDITS_NPH = 12,
  parameter        integer VC0_TOTAL_CREDITS_PD = 288,
  parameter        integer VC0_TOTAL_CREDITS_PH = 32,
  parameter        integer VC0_TX_LASTPACKET = 31,
  parameter [11:0] VC_BASE_PTR = 12'h10C,
  parameter [15:0] VC_CAP_ID = 16'h0002,
  parameter [11:0] VC_CAP_NEXTPTR = 12'h000,
  parameter        VC_CAP_ON = "FALSE",
  parameter        VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE",
  parameter [3:0]  VC_CAP_VERSION = 4'h1,
  parameter [11:0] VSEC_BASE_PTR = 12'h128,
  parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234,
  parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018,
  parameter [3:0]  VSEC_CAP_HDR_REVISION = 4'h1,
  parameter [15:0] VSEC_CAP_ID = 16'h000B,
  parameter        VSEC_CAP_IS_LINK_VISIBLE = "TRUE",
  parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140,
  parameter        VSEC_CAP_ON = "FALSE",
  parameter [3:0]  VSEC_CAP_VERSION = 4'h1
)
(
  input wire [C_DATA_WIDTH-1:0]         trn_td,
  input wire [REM_WIDTH-1:0]            trn_trem,
  input wire                trn_tsof,
  input wire                trn_teof,
  input wire                trn_tsrc_rdy,
  input wire                trn_tsrc_dsc,
  input wire                trn_terrfwd,
  input wire                trn_tecrc_gen,
  input wire                trn_tstr,
  input wire                trn_tcfg_gnt,
  input wire                trn_rdst_rdy,
  input wire                trn_rnp_req,
  input wire                trn_rfcp_ret,
  input wire                trn_rnp_ok,
  input wire        [2:0]   trn_fc_sel,
  input wire       [31:0]   trn_tdllp_data,
  input wire                trn_tdllp_src_rdy,
  input wire                ll2_tlp_rcv,
  input wire                ll2_send_enter_l1,
  input wire                ll2_send_enter_l23,
  input wire                ll2_send_as_req_l1,
  input wire                ll2_send_pm_ack,
  input wire        [4:0]   pl2_directed_lstate,
  input wire                ll2_suspend_now,
  input wire                tl2_ppm_suspend_req,
  input wire                tl2_aspm_suspend_credit_check,
  input wire        [1:0]   pl_directed_link_change,
  input wire        [1:0]   pl_directed_link_width,
  input wire                pl_directed_link_speed,
  input wire                pl_directed_link_auton,
  input wire                pl_upstream_prefer_deemph,
  input wire                pl_downstream_deemph_source,
  input wire                pl_directed_ltssm_new_vld,
  input wire        [5:0]   pl_directed_ltssm_new,
  input wire                pl_directed_ltssm_stall,
  input wire        [1:0]   pipe_rx0_char_is_k,
  input wire        [1:0]   pipe_rx1_char_is_k,
  input wire        [1:0]   pipe_rx2_char_is_k,
  input wire        [1:0]   pipe_rx3_char_is_k,
  input wire        [1:0]   pipe_rx4_char_is_k,
  input wire        [1:0]   pipe_rx5_char_is_k,
  input wire        [1:0]   pipe_rx6_char_is_k,
  input wire        [1:0]   pipe_rx7_char_is_k,
  input wire                pipe_rx0_valid,
  input wire                pipe_rx1_valid,
  input wire                pipe_rx2_valid,
  input wire                pipe_rx3_valid,
  input wire                pipe_rx4_valid,
  input wire                pipe_rx5_valid,
  input wire                pipe_rx6_valid,
  input wire                pipe_rx7_valid,
  input wire       [15:0]   pipe_rx0_data,
  input wire       [15:0]   pipe_rx1_data,
  input wire       [15:0]   pipe_rx2_data,
  input wire       [15:0]   pipe_rx3_data,
  input wire       [15:0]   pipe_rx4_data,
  input wire       [15:0]   pipe_rx5_data,
  input wire       [15:0]   pipe_rx6_data,
  input wire       [15:0]   pipe_rx7_data,
  input wire                pipe_rx0_chanisaligned,
  input wire                pipe_rx1_chanisaligned,
  input wire                pipe_rx2_chanisaligned,
  input wire                pipe_rx3_chanisaligned,
  input wire                pipe_rx4_chanisaligned,
  input wire                pipe_rx5_chanisaligned,
  input wire                pipe_rx6_chanisaligned,
  input wire                pipe_rx7_chanisaligned,
  input wire        [2:0]   pipe_rx0_status,
  input wire        [2:0]   pipe_rx1_status,
  input wire        [2:0]   pipe_rx2_status,
  input wire        [2:0]   pipe_rx3_status,
  input wire        [2:0]   pipe_rx4_status,
  input wire        [2:0]   pipe_rx5_status,
  input wire        [2:0]   pipe_rx6_status,
  input wire        [2:0]   pipe_rx7_status,
  input wire                pipe_rx0_phy_status,
  input wire                pipe_rx1_phy_status,
  input wire                pipe_rx2_phy_status,
  input wire                pipe_rx3_phy_status,
  input wire                pipe_rx4_phy_status,
  input wire                pipe_rx5_phy_status,
  input wire                pipe_rx6_phy_status,
  input wire                pipe_rx7_phy_status,
  input wire                pipe_rx0_elec_idle,
  input wire                pipe_rx1_elec_idle,
  input wire                pipe_rx2_elec_idle,
  input wire                pipe_rx3_elec_idle,
  input wire                pipe_rx4_elec_idle,
  input wire                pipe_rx5_elec_idle,
  input wire                pipe_rx6_elec_idle,
  input wire                pipe_rx7_elec_idle,
  input wire                pipe_clk,
  input wire                user_clk,
  input wire                user_clk2,
  input wire                user_clk_prebuf,
  input wire                user_clk_prebuf_en,
`ifdef B_TESTMODE
  input wire                scanmode_n,
  input wire                scanenable_n,
  input wire                edt_clk,
  input wire                edt_bypass,
  input wire                edt_update,
  input wire                edt_configuration,
  input wire                edt_single_bypass_chain,
  input wire                edt_channels_in1,
  input wire                edt_channels_in2,
  input wire                edt_channels_in3,
  input wire                edt_channels_in4,
  input wire                edt_channels_in5,
  input wire                edt_channels_in6,
  input wire                edt_channels_in7,
  input wire                edt_channels_in8,
  input wire                pmv_enable_n,
  input wire        [2:0]   pmv_select,
  input wire        [1:0]   pmv_divide,
`endif
  input wire                sys_rst_n,
  input wire                cm_rst_n,
  input wire                cm_sticky_rst_n,
  input wire                func_lvl_rst_n,
  input wire                tl_rst_n,
  input wire                dl_rst_n,
  input wire                pl_rst_n,
  input wire                pl_transmit_hot_rst,
//  input wire                cfg_reset,
//  input wire                gwe,
//  input wire                grestore,
//  input wire                ghigh,
  input wire       [31:0]   cfg_mgmt_di,
  input wire        [3:0]   cfg_mgmt_byte_en_n,
  input wire        [9:0]   cfg_mgmt_dwaddr,
  input wire                cfg_mgmt_wr_rw1c_as_rw_n,
  input wire                cfg_mgmt_wr_readonly_n,
  input wire                cfg_mgmt_wr_en_n,
  input wire                cfg_mgmt_rd_en_n,
  input wire                cfg_err_malformed_n,
  input wire                cfg_err_cor_n,
  input wire                cfg_err_ur_n,
  input wire                cfg_err_ecrc_n,
  input wire                cfg_err_cpl_timeout_n,
  input wire                cfg_err_cpl_abort_n,
  input wire                cfg_err_cpl_unexpect_n,
  input wire                cfg_err_poisoned_n,
  input wire                cfg_err_acs_n,
  input wire                cfg_err_atomic_egress_blocked_n,
  input wire                cfg_err_mc_blocked_n,
  input wire                cfg_err_internal_uncor_n,
  input wire                cfg_err_internal_cor_n,
  input wire                cfg_err_posted_n,
  input wire                cfg_err_locked_n,
  input wire                cfg_err_norecovery_n,
  input wire      [127:0]   cfg_err_aer_headerlog,
  input wire       [47:0]   cfg_err_tlp_cpl_header,
  input wire                cfg_interrupt_n,
  input wire        [7:0]   cfg_interrupt_di,
  input wire                cfg_interrupt_assert_n,
  input wire                cfg_interrupt_stat_n,
  input wire        [7:0]   cfg_ds_bus_number,
  input wire        [4:0]   cfg_ds_device_number,
  input wire        [2:0]   cfg_ds_function_number,
  input wire        [7:0]   cfg_port_number,
  input wire                cfg_pm_halt_aspm_l0s_n,
  input wire                cfg_pm_halt_aspm_l1_n,
  input wire                cfg_pm_force_state_en_n,
  input wire        [1:0]   cfg_pm_force_state,
  input wire                cfg_pm_wake_n,
  input wire                cfg_pm_turnoff_ok_n,
  input wire                cfg_pm_send_pme_to_n,
  input wire        [4:0]   cfg_pciecap_interrupt_msgnum,
  input wire                cfg_trn_pending_n,
  input wire        [2:0]   cfg_force_mps,
  input wire                cfg_force_common_clock_off,
  input wire                cfg_force_extended_sync_on,
  input wire       [63:0]   cfg_dsn,
  input wire        [4:0]   cfg_aer_interrupt_msgnum,
  input wire       [15:0]   cfg_dev_id,
  input wire       [15:0]   cfg_vend_id,
  input wire        [7:0]   cfg_rev_id,
  input wire       [15:0]   cfg_subsys_id,
  input wire       [15:0]   cfg_subsys_vend_id,
  input wire                drp_clk,
  input wire                drp_en,
  input wire                drp_we,
  input wire        [8:0]   drp_addr,
  input wire       [15:0]   drp_di,
  input wire        [1:0]   dbg_mode,
  input wire                dbg_sub_mode,
  input wire        [2:0]   pl_dbg_mode,

  output wire               trn_clk,

  output wire               trn_tdst_rdy,
  output wire               trn_terr_drop,
  output wire       [5:0]   trn_tbuf_av,
  output wire               trn_tcfg_req,

  //output wire [C_DATA_WIDTH-1:0]        trn_rd,
  output wire [127:0]        trn_rd,

  output wire [1:0]           trn_rrem,
  output wire               trn_rsof,
  output wire               trn_reof,
  output wire               trn_rsrc_rdy,
  output wire               trn_rsrc_dsc,
  output wire               trn_recrc_err,
  output wire               trn_rerrfwd,
  output wire       [7:0]   trn_rbar_hit,
  output wire               trn_lnk_up,
  output wire       [7:0]   trn_fc_ph,
  output wire      [11:0]   trn_fc_pd,
  output wire       [7:0]   trn_fc_nph,
  output wire      [11:0]   trn_fc_npd,
  output wire       [7:0]   trn_fc_cplh,
  output wire      [11:0]   trn_fc_cpld,
  output wire               trn_tdllp_dst_rdy,
  output wire      [63:0]   trn_rdllp_data,
  output wire       [1:0]   trn_rdllp_src_rdy,
  output wire               ll2_tfc_init1_seq,
  output wire               ll2_tfc_init2_seq,
  output wire               pl2_suspend_ok,
  output wire               pl2_recovery,
  output wire               pl2_rx_elec_idle,
  output wire       [1:0]   pl2_rx_pm_state,
  output wire               pl2_l0_req,
  output wire               ll2_suspend_ok,
  output wire               ll2_tx_idle,
  output wire       [4:0]   ll2_link_status,
  output wire               tl2_ppm_suspend_ok,
  output wire               tl2_aspm_suspend_req,
  output wire               tl2_aspm_suspend_credit_check_ok,
  output wire               pl2_link_up,
  output wire               pl2_receiver_err,
  output wire               ll2_receiver_err,
  output wire               ll2_protocol_err,
  output wire               ll2_bad_tlp_err,
  output wire               ll2_bad_dllp_err,
  output wire               ll2_replay_ro_err,
  output wire               ll2_replay_to_err,
  output wire      [63:0]   tl2_err_hdr,
  output wire               tl2_err_malformed,
  output wire               tl2_err_rxoverflow,
  output wire               tl2_err_fcpe,
  output wire               pl_sel_lnk_rate,
  output wire       [1:0]   pl_sel_lnk_width,
  output wire       [5:0]   pl_ltssm_state,
  output wire       [1:0]   pl_lane_reversal_mode,
  output wire               pl_phy_lnk_up_n,
  output wire       [2:0]   pl_tx_pm_state,
  output wire       [1:0]   pl_rx_pm_state,
  output wire               pl_link_upcfg_cap,
  output wire               pl_link_gen2_cap,
  output wire               pl_link_partner_gen2_supported,
  output wire       [2:0]   pl_initial_link_width,
  output wire               pl_directed_change_done,
  output wire               pipe_tx_rcvr_det,
  output wire               pipe_tx_reset,
  output wire               pipe_tx_rate,
  output wire               pipe_tx_deemph,
  output wire       [2:0]   pipe_tx_margin,
  output wire               pipe_rx0_polarity,
  output wire               pipe_rx1_polarity,
  output wire               pipe_rx2_polarity,
  output wire               pipe_rx3_polarity,
  output wire               pipe_rx4_polarity,
  output wire               pipe_rx5_polarity,
  output wire               pipe_rx6_polarity,
  output wire               pipe_rx7_polarity,
  output wire               pipe_tx0_compliance,
  output wire               pipe_tx1_compliance,
  output wire               pipe_tx2_compliance,
  output wire               pipe_tx3_compliance,
  output wire               pipe_tx4_compliance,
  output wire               pipe_tx5_compliance,
  output wire               pipe_tx6_compliance,
  output wire               pipe_tx7_compliance,
  output wire       [1:0]   pipe_tx0_char_is_k,
  output wire       [1:0]   pipe_tx1_char_is_k,
  output wire       [1:0]   pipe_tx2_char_is_k,
  output wire       [1:0]   pipe_tx3_char_is_k,
  output wire       [1:0]   pipe_tx4_char_is_k,
  output wire       [1:0]   pipe_tx5_char_is_k,
  output wire       [1:0]   pipe_tx6_char_is_k,
  output wire       [1:0]   pipe_tx7_char_is_k,
  output wire      [15:0]   pipe_tx0_data,
  output wire      [15:0]   pipe_tx1_data,
  output wire      [15:0]   pipe_tx2_data,
  output wire      [15:0]   pipe_tx3_data,
  output wire      [15:0]   pipe_tx4_data,
  output wire      [15:0]   pipe_tx5_data,
  output wire      [15:0]   pipe_tx6_data,
  output wire      [15:0]   pipe_tx7_data,
  output wire               pipe_tx0_elec_idle,
  output wire               pipe_tx1_elec_idle,
  output wire               pipe_tx2_elec_idle,
  output wire               pipe_tx3_elec_idle,
  output wire               pipe_tx4_elec_idle,
  output wire               pipe_tx5_elec_idle,
  output wire               pipe_tx6_elec_idle,
  output wire               pipe_tx7_elec_idle,
  output wire       [1:0]   pipe_tx0_powerdown,
  output wire       [1:0]   pipe_tx1_powerdown,
  output wire       [1:0]   pipe_tx2_powerdown,
  output wire       [1:0]   pipe_tx3_powerdown,
  output wire       [1:0]   pipe_tx4_powerdown,
  output wire       [1:0]   pipe_tx5_powerdown,
  output wire       [1:0]   pipe_tx6_powerdown,
  output wire       [1:0]   pipe_tx7_powerdown,
`ifdef B_TESTMODE
  output wire               pmv_out,
`endif
  output wire               user_rst_n,
  output wire               pl_received_hot_rst,
  output wire               received_func_lvl_rst_n,
  output wire               lnk_clk_en,
  output wire      [31:0]   cfg_mgmt_do,
  output wire               cfg_mgmt_rd_wr_done_n,
  output wire               cfg_err_aer_headerlog_set_n,
  output wire               cfg_err_cpl_rdy_n,
  output wire               cfg_interrupt_rdy_n,
  output wire       [2:0]   cfg_interrupt_mmenable,
  output wire               cfg_interrupt_msienable,
  output wire       [7:0]   cfg_interrupt_do,
  output wire               cfg_interrupt_msixenable,
  output wire               cfg_interrupt_msixfm,
  output wire               cfg_msg_received,
  output wire      [15:0]   cfg_msg_data,
  output wire               cfg_msg_received_err_cor,
  output wire               cfg_msg_received_err_non_fatal,
  output wire               cfg_msg_received_err_fatal,
  output wire               cfg_msg_received_assert_int_a,
  output wire               cfg_msg_received_deassert_int_a,
  output wire               cfg_msg_received_assert_int_b,
  output wire               cfg_msg_received_deassert_int_b,
  output wire               cfg_msg_received_assert_int_c,
  output wire               cfg_msg_received_deassert_int_c,
  output wire               cfg_msg_received_assert_int_d,
  output wire               cfg_msg_received_deassert_int_d,
  output wire               cfg_msg_received_pm_pme,
  output wire               cfg_msg_received_pme_to_ack,
  output wire               cfg_msg_received_pme_to,
  output wire               cfg_msg_received_setslotpowerlimit,
  output wire               cfg_msg_received_unlock,
  output wire               cfg_msg_received_pm_as_nak,
  output wire       [2:0]   cfg_pcie_link_state,
  output wire               cfg_pm_rcv_as_req_l1_n,
  output wire               cfg_pm_rcv_enter_l1_n,
  output wire               cfg_pm_rcv_enter_l23_n,
  output wire               cfg_pm_rcv_req_ack_n,
  output wire       [1:0]   cfg_pmcsr_powerstate,
  output wire               cfg_pmcsr_pme_en,
  output wire               cfg_pmcsr_pme_status,
  output wire               cfg_transaction,
  output wire               cfg_transaction_type,
  output wire       [6:0]   cfg_transaction_addr,
  output wire               cfg_command_io_enable,
  output wire               cfg_command_mem_enable,
  output wire               cfg_command_bus_master_enable,
  output wire               cfg_command_interrupt_disable,
  output wire               cfg_command_serr_en,
  output wire               cfg_bridge_serr_en,
  output wire               cfg_dev_status_corr_err_detected,
  output wire               cfg_dev_status_non_fatal_err_detected,
  output wire               cfg_dev_status_fatal_err_detected,
  output wire               cfg_dev_status_ur_detected,
  output wire               cfg_dev_control_corr_err_reporting_en,
  output wire               cfg_dev_control_non_fatal_reporting_en,
  output wire               cfg_dev_control_fatal_err_reporting_en,
  output wire               cfg_dev_control_ur_err_reporting_en,
  output wire               cfg_dev_control_enable_ro,
  output wire       [2:0]   cfg_dev_control_max_payload,
  output wire               cfg_dev_control_ext_tag_en,
  output wire               cfg_dev_control_phantom_en,
  output wire               cfg_dev_control_aux_power_en,
  output wire               cfg_dev_control_no_snoop_en,
  output wire       [2:0]   cfg_dev_control_max_read_req,
  output wire       [1:0]   cfg_link_status_current_speed,
  output wire       [3:0]   cfg_link_status_negotiated_width,
  output wire               cfg_link_status_link_training,
  output wire               cfg_link_status_dll_active,
  output wire               cfg_link_status_bandwidth_status,
  output wire               cfg_link_status_auto_bandwidth_status,
  output wire       [1:0]   cfg_link_control_aspm_control,
  output wire               cfg_link_control_rcb,
  output wire               cfg_link_control_link_disable,
  output wire               cfg_link_control_retrain_link,
  output wire               cfg_link_control_common_clock,
  output wire               cfg_link_control_extended_sync,
  output wire               cfg_link_control_clock_pm_en,
  output wire               cfg_link_control_hw_auto_width_dis,
  output wire               cfg_link_control_bandwidth_int_en,
  output wire               cfg_link_control_auto_bandwidth_int_en,
  output wire       [3:0]   cfg_dev_control2_cpl_timeout_val,
  output wire               cfg_dev_control2_cpl_timeout_dis,
  output wire               cfg_dev_control2_ari_forward_en,
  output wire               cfg_dev_control2_atomic_requester_en,
  output wire               cfg_dev_control2_atomic_egress_block,
  output wire               cfg_dev_control2_ido_req_en,
  output wire               cfg_dev_control2_ido_cpl_en,
  output wire               cfg_dev_control2_ltr_en,
  output wire               cfg_dev_control2_tlp_prefix_block,
  output wire               cfg_slot_control_electromech_il_ctl_pulse,
  output wire               cfg_root_control_syserr_corr_err_en,
  output wire               cfg_root_control_syserr_non_fatal_err_en,
  output wire               cfg_root_control_syserr_fatal_err_en,
  output wire               cfg_root_control_pme_int_en,
  output wire               cfg_aer_ecrc_check_en,
  output wire               cfg_aer_ecrc_gen_en,
  output wire               cfg_aer_rooterr_corr_err_reporting_en,
  output wire               cfg_aer_rooterr_non_fatal_err_reporting_en,
  output wire               cfg_aer_rooterr_fatal_err_reporting_en,
  output wire               cfg_aer_rooterr_corr_err_received,
  output wire               cfg_aer_rooterr_non_fatal_err_received,
  output wire               cfg_aer_rooterr_fatal_err_received,
  output wire       [6:0]   cfg_vc_tcvc_map,
  output wire               drp_rdy,
  output wire      [15:0]   drp_do,
  output wire      [63:0]   dbg_vec_a,
  output wire      [63:0]   dbg_vec_b,
  output wire      [11:0]   dbg_vec_c,
  output wire               dbg_sclr_a,
  output wire               dbg_sclr_b,
  output wire               dbg_sclr_c,
  output wire               dbg_sclr_d,
  output wire               dbg_sclr_e,
  output wire               dbg_sclr_f,
  output wire               dbg_sclr_g,
  output wire               dbg_sclr_h,
  output wire               dbg_sclr_i,
  output wire               dbg_sclr_j,
  output wire               dbg_sclr_k,
  output wire      [11:0]   pl_dbg_vec
//  output wire      [18:0]   xil_unconn_out
);

  localparam        TCQ = 1;

  wire [3:0]        trn_tdst_rdy_bus;

  // Assignments to outputs
  assign            trn_clk = user_clk2;
  assign            trn_tdst_rdy = trn_tdst_rdy_bus[0];

  //----------------------------------------------------------------------//
  // BRAM                                                                 //
  //----------------------------------------------------------------------//

  // transmit bram interface
  wire        mim_tx_wen;
  wire [12:0] mim_tx_waddr;
  wire [68:0] mim_tx_wdata;
  wire        mim_tx_ren;
  wire        mim_tx_rce;
  wire [12:0] mim_tx_raddr;
  wire [68:0] mim_tx_rdata;
  wire [2:0]  unused_mim_tx_rdata;

  // receive bram interface
  wire        mim_rx_wen;
  wire [12:0] mim_rx_waddr;
  wire [67:0] mim_rx_wdata;
  wire        mim_rx_ren;
  wire        mim_rx_rce;
  wire [12:0] mim_rx_raddr;
  wire [67:0] mim_rx_rdata;
  wire [3:0]  unused_mim_rx_rdata;

model_ap2_tst_pcie_bram_top_7x #(
    .LINK_CAP_MAX_LINK_SPEED       ( LINK_CAP_MAX_LINK_SPEED ),
    .LINK_CAP_MAX_LINK_WIDTH       ( LINK_CAP_MAX_LINK_WIDTH ),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED ( DEV_CAP_MAX_PAYLOAD_SUPPORTED ),
    .VC0_TX_LASTPACKET             ( VC0_TX_LASTPACKET ),
    .TL_TX_RAM_RADDR_LATENCY       ( TL_TX_RAM_RADDR_LATENCY ),
    .TL_TX_RAM_RDATA_LATENCY       ( TL_TX_RAM_RDATA_LATENCY ),
    .TL_TX_RAM_WRITE_LATENCY       ( TL_TX_RAM_WRITE_LATENCY ),
    .VC0_RX_RAM_LIMIT              ( VC0_RX_RAM_LIMIT ),
    .TL_RX_RAM_RADDR_LATENCY       ( TL_RX_RAM_RADDR_LATENCY ),
    .TL_RX_RAM_RDATA_LATENCY       ( TL_RX_RAM_RDATA_LATENCY ),
    .TL_RX_RAM_WRITE_LATENCY       ( TL_RX_RAM_WRITE_LATENCY )
  ) model_ap2_tst_pcie_bram_top (
    .user_clk_i    ( user_clk ),
    .reset_i       ( 1'b0 ),

    .mim_tx_waddr  ( mim_tx_waddr ),
    .mim_tx_wen    ( mim_tx_wen ),
    .mim_tx_ren    ( mim_tx_ren ),
    .mim_tx_rce    ( 1'b1 ),
    .mim_tx_wdata  ( {3'b0, mim_tx_wdata} ),
    .mim_tx_raddr  ( mim_tx_raddr ),
    .mim_tx_rdata  ( {unused_mim_tx_rdata, mim_tx_rdata} ),

    .mim_rx_waddr  ( mim_rx_waddr ),
    .mim_rx_wen    ( mim_rx_wen ),
    .mim_rx_ren    ( mim_rx_ren ),
    .mim_rx_rce    ( 1'b1 ),
    .mim_rx_wdata  ( {4'b0, mim_rx_wdata} ),
    .mim_rx_raddr  ( mim_rx_raddr ),
    .mim_rx_rdata  ( {unused_mim_rx_rdata, mim_rx_rdata} )
 );

  //-------------------------------------------------------
  // Virtex7 PCI Express Block Module
  //-------------------------------------------------------

  PCIE_2_1 #(  // Verilog-2001
    .AER_BASE_PTR                             ( AER_BASE_PTR ),
    .AER_CAP_ECRC_CHECK_CAPABLE               ( AER_CAP_ECRC_CHECK_CAPABLE ),
    .AER_CAP_ECRC_GEN_CAPABLE                 ( AER_CAP_ECRC_GEN_CAPABLE ),
    .AER_CAP_ID                               ( AER_CAP_ID ),
    .AER_CAP_MULTIHEADER                      ( AER_CAP_MULTIHEADER ),
    .AER_CAP_NEXTPTR                          ( AER_CAP_NEXTPTR ),
    .AER_CAP_ON                               ( AER_CAP_ON ),
    .AER_CAP_OPTIONAL_ERR_SUPPORT             ( AER_CAP_OPTIONAL_ERR_SUPPORT ),
    .AER_CAP_PERMIT_ROOTERR_UPDATE            ( AER_CAP_PERMIT_ROOTERR_UPDATE ),
    .AER_CAP_VERSION                          ( AER_CAP_VERSION ),
    .ALLOW_X8_GEN2                            ( ALLOW_X8_GEN2 ),
    .BAR0                                     ( BAR0 ),
    .BAR1                                     ( BAR1 ),
    .BAR2                                     ( BAR2 ),
    .BAR3                                     ( BAR3 ),
    .BAR4                                     ( BAR4 ),
    .BAR5                                     ( BAR5 ),
    .CAPABILITIES_PTR                         ( CAPABILITIES_PTR ),
    .CARDBUS_CIS_POINTER                      ( CARDBUS_CIS_POINTER ),
    .CFG_ECRC_ERR_CPLSTAT                     ( CFG_ECRC_ERR_CPLSTAT ),
    .CLASS_CODE                               ( CLASS_CODE ),
    .CMD_INTX_IMPLEMENTED                     ( CMD_INTX_IMPLEMENTED ),
    .CPL_TIMEOUT_DISABLE_SUPPORTED            ( CPL_TIMEOUT_DISABLE_SUPPORTED ),
    .CPL_TIMEOUT_RANGES_SUPPORTED             ( CPL_TIMEOUT_RANGES_SUPPORTED ),
    .CRM_MODULE_RSTS                          ( CRM_MODULE_RSTS ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE ),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      ( DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE ),
    .DEV_CAP_ENDPOINT_L0S_LATENCY             ( DEV_CAP_ENDPOINT_L0S_LATENCY ),
    .DEV_CAP_ENDPOINT_L1_LATENCY              ( DEV_CAP_ENDPOINT_L1_LATENCY ),
    .DEV_CAP_EXT_TAG_SUPPORTED                ( DEV_CAP_EXT_TAG_SUPPORTED ),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     ( DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE ),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED            ( DEV_CAP_MAX_PAYLOAD_SUPPORTED ),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        ( DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT ),
    .DEV_CAP_ROLE_BASED_ERROR                 ( DEV_CAP_ROLE_BASED_ERROR ),
    .DEV_CAP_RSVD_14_12                       ( DEV_CAP_RSVD_14_12 ),
    .DEV_CAP_RSVD_17_16                       ( DEV_CAP_RSVD_17_16 ),
    .DEV_CAP_RSVD_31_29                       ( DEV_CAP_RSVD_31_29 ),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED        ( DEV_CAP2_ARI_FORWARDING_SUPPORTED ),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      ( DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED ),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  ( DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED ),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED      ( DEV_CAP2_CAS128_COMPLETER_SUPPORTED ),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     ( DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED ),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    ( DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED ),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED         ( DEV_CAP2_LTR_MECHANISM_SUPPORTED ),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         ( DEV_CAP2_MAX_ENDEND_TLP_PREFIXES ),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      ( DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING ),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED         ( DEV_CAP2_TPH_COMPLETER_SUPPORTED ),
    .DEV_CONTROL_AUX_POWER_SUPPORTED          ( DEV_CONTROL_AUX_POWER_SUPPORTED ),
    .DEV_CONTROL_EXT_TAG_DEFAULT              ( DEV_CONTROL_EXT_TAG_DEFAULT ),
    .DISABLE_ASPM_L1_TIMER                    ( DISABLE_ASPM_L1_TIMER ),
    .DISABLE_BAR_FILTERING                    ( DISABLE_BAR_FILTERING ),
    .DISABLE_ERR_MSG                          ( DISABLE_ERR_MSG ),
    .DISABLE_ID_CHECK                         ( DISABLE_ID_CHECK ),
    .DISABLE_LANE_REVERSAL                    ( DISABLE_LANE_REVERSAL ),
    .DISABLE_LOCKED_FILTER                    ( DISABLE_LOCKED_FILTER ),
    .DISABLE_PPM_FILTER                       ( DISABLE_PPM_FILTER ),
    .DISABLE_RX_POISONED_RESP                 ( DISABLE_RX_POISONED_RESP ),
    .DISABLE_RX_TC_FILTER                     ( DISABLE_RX_TC_FILTER ),
    .DISABLE_SCRAMBLING                       ( DISABLE_SCRAMBLING ),
    .DNSTREAM_LINK_NUM                        ( DNSTREAM_LINK_NUM ),
    .DSN_BASE_PTR                             ( DSN_BASE_PTR ),
    .DSN_CAP_ID                               ( DSN_CAP_ID ),
    .DSN_CAP_NEXTPTR                          ( DSN_CAP_NEXTPTR ),
    .DSN_CAP_ON                               ( DSN_CAP_ON ),
    .DSN_CAP_VERSION                          ( DSN_CAP_VERSION ),
    .ENABLE_MSG_ROUTE                         ( ENABLE_MSG_ROUTE ),
    .ENABLE_RX_TD_ECRC_TRIM                   ( ENABLE_RX_TD_ECRC_TRIM ),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   ( ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED ),
    .ENTER_RVRY_EI_L0                         ( ENTER_RVRY_EI_L0 ),
    .EXIT_LOOPBACK_ON_EI                      ( EXIT_LOOPBACK_ON_EI ),
    .EXPANSION_ROM                            ( EXPANSION_ROM ),
    .EXT_CFG_CAP_PTR                          ( EXT_CFG_CAP_PTR ),
    .EXT_CFG_XP_CAP_PTR                       ( EXT_CFG_XP_CAP_PTR ),
    .HEADER_TYPE                              ( HEADER_TYPE ),
    .INFER_EI                                 ( INFER_EI ),
    .INTERRUPT_PIN                            ( INTERRUPT_PIN ),
    .INTERRUPT_STAT_AUTO                      ( INTERRUPT_STAT_AUTO ),
    .IS_SWITCH                                ( IS_SWITCH ),
    .LAST_CONFIG_DWORD                        ( LAST_CONFIG_DWORD ),
    .LINK_CAP_ASPM_OPTIONALITY                ( LINK_CAP_ASPM_OPTIONALITY ),
    .LINK_CAP_ASPM_SUPPORT                    ( LINK_CAP_ASPM_SUPPORT ),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT          ( LINK_CAP_CLOCK_POWER_MANAGEMENT ),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   ( LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP ),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ( LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    ( LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1           ( LINK_CAP_L0S_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2           ( LINK_CAP_L0S_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     ( LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1            ( LINK_CAP_L1_EXIT_LATENCY_GEN1 ),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2            ( LINK_CAP_L1_EXIT_LATENCY_GEN2 ),
    .LINK_CAP_MAX_LINK_SPEED                  ( LINK_CAP_MAX_LINK_SPEED ),
    .LINK_CAP_MAX_LINK_WIDTH                  ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_RSVD_23                         ( LINK_CAP_RSVD_23 ),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     ( LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE ),
    .LINK_CONTROL_RCB                         ( LINK_CONTROL_RCB ),
    .LINK_CTRL2_DEEMPHASIS                    ( LINK_CTRL2_DEEMPHASIS ),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   ( LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE ),
    .LINK_CTRL2_TARGET_LINK_SPEED             ( LINK_CTRL2_TARGET_LINK_SPEED ),
    .LINK_STATUS_SLOT_CLOCK_CONFIG            ( LINK_STATUS_SLOT_CLOCK_CONFIG ),
    .LL_ACK_TIMEOUT                           ( LL_ACK_TIMEOUT ),
    .LL_ACK_TIMEOUT_EN                        ( LL_ACK_TIMEOUT_EN ),
    .LL_ACK_TIMEOUT_FUNC                      ( LL_ACK_TIMEOUT_FUNC ),
    .LL_REPLAY_TIMEOUT                        ( LL_REPLAY_TIMEOUT ),
    .LL_REPLAY_TIMEOUT_EN                     ( LL_REPLAY_TIMEOUT_EN ),
    .LL_REPLAY_TIMEOUT_FUNC                   ( LL_REPLAY_TIMEOUT_FUNC ),
    .LTSSM_MAX_LINK_WIDTH                     ( LTSSM_MAX_LINK_WIDTH ),
    .MPS_FORCE                                ( MPS_FORCE ),
    .MSI_BASE_PTR                             ( MSI_BASE_PTR ),
    .MSI_CAP_ID                               ( MSI_CAP_ID ),
    .MSI_CAP_MULTIMSG_EXTENSION               ( MSI_CAP_MULTIMSG_EXTENSION ),
    .MSI_CAP_MULTIMSGCAP                      ( MSI_CAP_MULTIMSGCAP ),
    .MSI_CAP_NEXTPTR                          ( MSI_CAP_NEXTPTR ),
    .MSI_CAP_ON                               ( MSI_CAP_ON ),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE       ( MSI_CAP_PER_VECTOR_MASKING_CAPABLE ),
    .MSI_CAP_64_BIT_ADDR_CAPABLE              ( MSI_CAP_64_BIT_ADDR_CAPABLE ),
    .MSIX_BASE_PTR                            ( MSIX_BASE_PTR ),
    .MSIX_CAP_ID                              ( MSIX_CAP_ID ),
    .MSIX_CAP_NEXTPTR                         ( MSIX_CAP_NEXTPTR ),
    .MSIX_CAP_ON                              ( MSIX_CAP_ON ),
    .MSIX_CAP_PBA_BIR                         ( MSIX_CAP_PBA_BIR ),
    .MSIX_CAP_PBA_OFFSET                      ( MSIX_CAP_PBA_OFFSET ),
    .MSIX_CAP_TABLE_BIR                       ( MSIX_CAP_TABLE_BIR ),
    .MSIX_CAP_TABLE_OFFSET                    ( MSIX_CAP_TABLE_OFFSET ),
    .MSIX_CAP_TABLE_SIZE                      ( MSIX_CAP_TABLE_SIZE ),
    .N_FTS_COMCLK_GEN1                        ( N_FTS_COMCLK_GEN1 ),
    .N_FTS_COMCLK_GEN2                        ( N_FTS_COMCLK_GEN2 ),
    .N_FTS_GEN1                               ( N_FTS_GEN1 ),
    .N_FTS_GEN2                               ( N_FTS_GEN2 ),
    .PCIE_BASE_PTR                            ( PCIE_BASE_PTR ),
    .PCIE_CAP_CAPABILITY_ID                   ( PCIE_CAP_CAPABILITY_ID ),
    .PCIE_CAP_CAPABILITY_VERSION              ( PCIE_CAP_CAPABILITY_VERSION ),
    .PCIE_CAP_DEVICE_PORT_TYPE                ( PCIE_CAP_DEVICE_PORT_TYPE ),
    .PCIE_CAP_NEXTPTR                         ( PCIE_CAP_NEXTPTR ),
    .PCIE_CAP_ON                              ( PCIE_CAP_ON ),
    .PCIE_CAP_RSVD_15_14                      ( PCIE_CAP_RSVD_15_14 ),
    .PCIE_CAP_SLOT_IMPLEMENTED                ( PCIE_CAP_SLOT_IMPLEMENTED ),
    .PCIE_REVISION                            ( PCIE_REVISION ),
    .PL_AUTO_CONFIG                           ( PL_AUTO_CONFIG ),
    .PL_FAST_TRAIN                            ( PL_FAST_TRAIN ),
    .PM_ASPML0S_TIMEOUT                       ( PM_ASPML0S_TIMEOUT ),
    .PM_ASPML0S_TIMEOUT_EN                    ( PM_ASPML0S_TIMEOUT_EN ),
    .PM_ASPML0S_TIMEOUT_FUNC                  ( PM_ASPML0S_TIMEOUT_FUNC ),
    .PM_ASPM_FASTEXIT                         ( PM_ASPM_FASTEXIT ),
    .PM_BASE_PTR                              ( PM_BASE_PTR ),
    .PM_CAP_AUXCURRENT                        ( PM_CAP_AUXCURRENT ),
    .PM_CAP_DSI                               ( PM_CAP_DSI ),
    .PM_CAP_D1SUPPORT                         ( PM_CAP_D1SUPPORT ),
    .PM_CAP_D2SUPPORT                         ( PM_CAP_D2SUPPORT ),
    .PM_CAP_ID                                ( PM_CAP_ID ),
    .PM_CAP_NEXTPTR                           ( PM_CAP_NEXTPTR ),
    .PM_CAP_ON                                ( PM_CAP_ON ),
    .PM_CAP_PME_CLOCK                         ( PM_CAP_PME_CLOCK ),
    .PM_CAP_PMESUPPORT                        ( PM_CAP_PMESUPPORT ),
    .PM_CAP_RSVD_04                           ( PM_CAP_RSVD_04 ),
    .PM_CAP_VERSION                           ( PM_CAP_VERSION ),
    .PM_CSR_BPCCEN                            ( PM_CSR_BPCCEN ),
    .PM_CSR_B2B3                              ( PM_CSR_B2B3 ),
    .PM_CSR_NOSOFTRST                         ( PM_CSR_NOSOFTRST ),
    .PM_DATA_SCALE0                           ( PM_DATA_SCALE0 ),
    .PM_DATA_SCALE1                           ( PM_DATA_SCALE1 ),
    .PM_DATA_SCALE2                           ( PM_DATA_SCALE2 ),
    .PM_DATA_SCALE3                           ( PM_DATA_SCALE3 ),
    .PM_DATA_SCALE4                           ( PM_DATA_SCALE4 ),
    .PM_DATA_SCALE5                           ( PM_DATA_SCALE5 ),
    .PM_DATA_SCALE6                           ( PM_DATA_SCALE6 ),
    .PM_DATA_SCALE7                           ( PM_DATA_SCALE7 ),
    .PM_DATA0                                 ( PM_DATA0 ),
    .PM_DATA1                                 ( PM_DATA1 ),
    .PM_DATA2                                 ( PM_DATA2 ),
    .PM_DATA3                                 ( PM_DATA3 ),
    .PM_DATA4                                 ( PM_DATA4 ),
    .PM_DATA5                                 ( PM_DATA5 ),
    .PM_DATA6                                 ( PM_DATA6 ),
    .PM_DATA7                                 ( PM_DATA7 ),
    .PM_MF                                    ( PM_MF ),
    .RBAR_BASE_PTR                            ( RBAR_BASE_PTR ),
    .RBAR_CAP_CONTROL_ENCODEDBAR0             ( RBAR_CAP_CONTROL_ENCODEDBAR0 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR1             ( RBAR_CAP_CONTROL_ENCODEDBAR1 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR2             ( RBAR_CAP_CONTROL_ENCODEDBAR2 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR3             ( RBAR_CAP_CONTROL_ENCODEDBAR3 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR4             ( RBAR_CAP_CONTROL_ENCODEDBAR4 ),
    .RBAR_CAP_CONTROL_ENCODEDBAR5             ( RBAR_CAP_CONTROL_ENCODEDBAR5 ),
    .RBAR_CAP_ID                              ( RBAR_CAP_ID ),
    .RBAR_CAP_INDEX0                          ( RBAR_CAP_INDEX0 ),
    .RBAR_CAP_INDEX1                          ( RBAR_CAP_INDEX1 ),
    .RBAR_CAP_INDEX2                          ( RBAR_CAP_INDEX2 ),
    .RBAR_CAP_INDEX3                          ( RBAR_CAP_INDEX3 ),
    .RBAR_CAP_INDEX4                          ( RBAR_CAP_INDEX4 ),
    .RBAR_CAP_INDEX5                          ( RBAR_CAP_INDEX5 ),
    .RBAR_CAP_NEXTPTR                         ( RBAR_CAP_NEXTPTR ),
    .RBAR_CAP_ON                              ( RBAR_CAP_ON ),
    .RBAR_CAP_SUP0                            ( RBAR_CAP_SUP0 ),
    .RBAR_CAP_SUP1                            ( RBAR_CAP_SUP1 ),
    .RBAR_CAP_SUP2                            ( RBAR_CAP_SUP2 ),
    .RBAR_CAP_SUP3                            ( RBAR_CAP_SUP3 ),
    .RBAR_CAP_SUP4                            ( RBAR_CAP_SUP4 ),
    .RBAR_CAP_SUP5                            ( RBAR_CAP_SUP5 ),
    .RBAR_CAP_VERSION                         ( RBAR_CAP_VERSION ),
    .RBAR_NUM                                 ( RBAR_NUM ),
    .RECRC_CHK                                ( RECRC_CHK ),
    .RECRC_CHK_TRIM                           ( RECRC_CHK_TRIM ),
    .ROOT_CAP_CRS_SW_VISIBILITY               ( ROOT_CAP_CRS_SW_VISIBILITY ),
    .RP_AUTO_SPD                              ( RP_AUTO_SPD ),
    .RP_AUTO_SPD_LOOPCNT                      ( RP_AUTO_SPD_LOOPCNT ),
    .SELECT_DLL_IF                            ( SELECT_DLL_IF ),
    .SLOT_CAP_ATT_BUTTON_PRESENT              ( SLOT_CAP_ATT_BUTTON_PRESENT ),
    .SLOT_CAP_ATT_INDICATOR_PRESENT           ( SLOT_CAP_ATT_INDICATOR_PRESENT ),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT          ( SLOT_CAP_ELEC_INTERLOCK_PRESENT ),
    .SLOT_CAP_HOTPLUG_CAPABLE                 ( SLOT_CAP_HOTPLUG_CAPABLE ),
    .SLOT_CAP_HOTPLUG_SURPRISE                ( SLOT_CAP_HOTPLUG_SURPRISE ),
    .SLOT_CAP_MRL_SENSOR_PRESENT              ( SLOT_CAP_MRL_SENSOR_PRESENT ),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        ( SLOT_CAP_NO_CMD_COMPLETED_SUPPORT ),
    .SLOT_CAP_PHYSICAL_SLOT_NUM               ( SLOT_CAP_PHYSICAL_SLOT_NUM ),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT        ( SLOT_CAP_POWER_CONTROLLER_PRESENT ),
    .SLOT_CAP_POWER_INDICATOR_PRESENT         ( SLOT_CAP_POWER_INDICATOR_PRESENT ),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE          ( SLOT_CAP_SLOT_POWER_LIMIT_SCALE ),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE          ( SLOT_CAP_SLOT_POWER_LIMIT_VALUE ),
    .SPARE_BIT0                               ( SPARE_BIT0 ),
    .SPARE_BIT1                               ( SPARE_BIT1 ),
    .SPARE_BIT2                               ( SPARE_BIT2 ),
    .SPARE_BIT3                               ( SPARE_BIT3 ),
    .SPARE_BIT4                               ( SPARE_BIT4 ),
    .SPARE_BIT5                               ( SPARE_BIT5 ),
    .SPARE_BIT6                               ( SPARE_BIT6 ),
    .SPARE_BIT7                               ( SPARE_BIT7 ),
    .SPARE_BIT8                               ( SPARE_BIT8 ),
    .SPARE_BYTE0                              ( SPARE_BYTE0 ),
    .SPARE_BYTE1                              ( SPARE_BYTE1 ),
    .SPARE_BYTE2                              ( SPARE_BYTE2 ),
    .SPARE_BYTE3                              ( SPARE_BYTE3 ),
    .SPARE_WORD0                              ( SPARE_WORD0 ),
    .SPARE_WORD1                              ( SPARE_WORD1 ),
    .SPARE_WORD2                              ( SPARE_WORD2 ),
    .SPARE_WORD3                              ( SPARE_WORD3 ),
    .SSL_MESSAGE_AUTO                         ( SSL_MESSAGE_AUTO ),
    .TECRC_EP_INV                             ( TECRC_EP_INV ),
    .TL_RBYPASS                               ( TL_RBYPASS ),
    .TL_RX_RAM_RADDR_LATENCY                  ( TL_RX_RAM_RADDR_LATENCY ),
    .TL_RX_RAM_RDATA_LATENCY                  ( TL_RX_RAM_RDATA_LATENCY ),
    .TL_RX_RAM_WRITE_LATENCY                  ( TL_RX_RAM_WRITE_LATENCY ),
    .TL_TFC_DISABLE                           ( TL_TFC_DISABLE ),
    .TL_TX_CHECKS_DISABLE                     ( TL_TX_CHECKS_DISABLE ),
    .TL_TX_RAM_RADDR_LATENCY                  ( TL_TX_RAM_RADDR_LATENCY ),
    .TL_TX_RAM_RDATA_LATENCY                  ( TL_TX_RAM_RDATA_LATENCY ),
    .TL_TX_RAM_WRITE_LATENCY                  ( TL_TX_RAM_WRITE_LATENCY ),
    .TRN_DW                                   ( TRN_DW ),
    .TRN_NP_FC                                ( TRN_NP_FC ),
    .UPCONFIG_CAPABLE                         ( UPCONFIG_CAPABLE ),
    .UPSTREAM_FACING                          ( UPSTREAM_FACING ),
    .UR_ATOMIC                                ( UR_ATOMIC ),
    .UR_CFG1                                  ( UR_CFG1 ),
    .UR_INV_REQ                               ( UR_INV_REQ ),
    .UR_PRS_RESPONSE                          ( UR_PRS_RESPONSE ),
    .USE_RID_PINS                             ( USE_RID_PINS ),
    .USER_CLK_FREQ                            ( USER_CLK_FREQ ),
    .USER_CLK2_DIV2                           ( USER_CLK2_DIV2 ),
    .VC_BASE_PTR                              ( VC_BASE_PTR ),
    .VC_CAP_ID                                ( VC_CAP_ID ),
    .VC_CAP_NEXTPTR                           ( VC_CAP_NEXTPTR ),
    .VC_CAP_ON                                ( VC_CAP_ON ),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS         ( VC_CAP_REJECT_SNOOP_TRANSACTIONS ),
    .VC_CAP_VERSION                           ( VC_CAP_VERSION ),
    .VC0_CPL_INFINITE                         ( VC0_CPL_INFINITE ),
    .VC0_RX_RAM_LIMIT                         ( VC0_RX_RAM_LIMIT ),
    .VC0_TOTAL_CREDITS_CD                     ( VC0_TOTAL_CREDITS_CD ),
    .VC0_TOTAL_CREDITS_CH                     ( VC0_TOTAL_CREDITS_CH ),
    .VC0_TOTAL_CREDITS_NPD                    ( VC0_TOTAL_CREDITS_NPD ),
    .VC0_TOTAL_CREDITS_NPH                    ( VC0_TOTAL_CREDITS_NPH ),
    .VC0_TOTAL_CREDITS_PD                     ( VC0_TOTAL_CREDITS_PD ),
    .VC0_TOTAL_CREDITS_PH                     ( VC0_TOTAL_CREDITS_PH ),
    .VC0_TX_LASTPACKET                        ( VC0_TX_LASTPACKET ),
    .VSEC_BASE_PTR                            ( VSEC_BASE_PTR ),
    .VSEC_CAP_HDR_ID                          ( VSEC_CAP_HDR_ID ),
    .VSEC_CAP_HDR_REVISION                    ( VSEC_CAP_HDR_REVISION ),
    .VSEC_CAP_ID                              ( VSEC_CAP_ID ),
    .VSEC_CAP_IS_LINK_VISIBLE                 ( VSEC_CAP_IS_LINK_VISIBLE ),
    .VSEC_CAP_NEXTPTR                         ( VSEC_CAP_NEXTPTR ),
    .VSEC_CAP_ON                              ( VSEC_CAP_ON ),
    .VSEC_CAP_VERSION                         ( VSEC_CAP_VERSION )
`ifdef B_TESTMODE
    ,
    .TEST_MODE_PIN_CHAR                       ( TEST_MODE_PIN_CHAR )
`endif

  )
  pcie_block_i (
  
    .TRNTD                               (trn_td                                     ),
    .TRNTREM                             (trn_trem                                   ),


    .TRNTSOF                             (trn_tsof                                   ),
    .TRNTEOF                             (trn_teof                                   ),
    .TRNTSRCRDY                          (trn_tsrc_rdy                               ),
    .TRNTSRCDSC                          (trn_tsrc_dsc                               ),
    .TRNTERRFWD                          (trn_terrfwd                                ),
    .TRNTECRCGEN                         (trn_tecrc_gen                              ),
    .TRNTSTR                             (trn_tstr                                   ),
    .TRNTCFGGNT                          (trn_tcfg_gnt                               ),
    .TRNRDSTRDY                          (trn_rdst_rdy                               ),
    .TRNRNPREQ                           (trn_rnp_req                                ),
    .TRNRFCPRET                          (trn_rfcp_ret                               ),
    .TRNRNPOK                            (trn_rnp_ok                                 ),
    .TRNFCSEL                            (trn_fc_sel                                 ),
    .MIMTXRDATA                          (mim_tx_rdata                               ),
    .MIMRXRDATA                          (mim_rx_rdata                               ),
    .TRNTDLLPDATA                        (trn_tdllp_data                             ),
    .TRNTDLLPSRCRDY                      (trn_tdllp_src_rdy                          ),
    .LL2TLPRCV                           (ll2_tlp_rcv                                ),
    .LL2SENDENTERL1                      (ll2_send_enter_l1                          ),
    .LL2SENDENTERL23                     (ll2_send_enter_l23                         ),
    .LL2SENDASREQL1                      (ll2_send_as_req_l1                         ),
    .LL2SENDPMACK                        (ll2_send_pm_ack                            ),
    .PL2DIRECTEDLSTATE                   (pl2_directed_lstate                        ),
    .LL2SUSPENDNOW                       (ll2_suspend_now                            ),
    .TL2PPMSUSPENDREQ                    (tl2_ppm_suspend_req                        ),
    .TL2ASPMSUSPENDCREDITCHECK           (tl2_aspm_suspend_credit_check              ),
    .PLDIRECTEDLINKCHANGE                (pl_directed_link_change                    ),
    .PLDIRECTEDLINKWIDTH                 (pl_directed_link_width                     ),
    .PLDIRECTEDLINKSPEED                 (pl_directed_link_speed                     ),
    .PLDIRECTEDLINKAUTON                 (pl_directed_link_auton                     ),
    .PLUPSTREAMPREFERDEEMPH              (pl_upstream_prefer_deemph                  ),
    .PLDOWNSTREAMDEEMPHSOURCE            (pl_downstream_deemph_source                ),
    .PLDIRECTEDLTSSMNEW                  (pl_directed_ltssm_new                      ),
    .PLDIRECTEDLTSSMNEWVLD               (pl_directed_ltssm_new_vld                  ),
    .PLDIRECTEDLTSSMSTALL                (pl_directed_ltssm_stall                    ),
    .PIPERX0CHARISK                      (pipe_rx0_char_is_k                         ),
    .PIPERX1CHARISK                      (pipe_rx1_char_is_k                         ),
    .PIPERX2CHARISK                      (pipe_rx2_char_is_k                         ),
    .PIPERX3CHARISK                      (pipe_rx3_char_is_k                         ),
    .PIPERX4CHARISK                      (pipe_rx4_char_is_k                         ),
    .PIPERX5CHARISK                      (pipe_rx5_char_is_k                         ),
    .PIPERX6CHARISK                      (pipe_rx6_char_is_k                         ),
    .PIPERX7CHARISK                      (pipe_rx7_char_is_k                         ),
    .PIPERX0VALID                        (pipe_rx0_valid                             ),
    .PIPERX1VALID                        (pipe_rx1_valid                             ),
    .PIPERX2VALID                        (pipe_rx2_valid                             ),
    .PIPERX3VALID                        (pipe_rx3_valid                             ),
    .PIPERX4VALID                        (pipe_rx4_valid                             ),
    .PIPERX5VALID                        (pipe_rx5_valid                             ),
    .PIPERX6VALID                        (pipe_rx6_valid                             ),
    .PIPERX7VALID                        (pipe_rx7_valid                             ),
    .PIPERX0DATA                         (pipe_rx0_data                              ),
    .PIPERX1DATA                         (pipe_rx1_data                              ),
    .PIPERX2DATA                         (pipe_rx2_data                              ),
    .PIPERX3DATA                         (pipe_rx3_data                              ),
    .PIPERX4DATA                         (pipe_rx4_data                              ),
    .PIPERX5DATA                         (pipe_rx5_data                              ),
    .PIPERX6DATA                         (pipe_rx6_data                              ),
    .PIPERX7DATA                         (pipe_rx7_data                              ),
    .PIPERX0CHANISALIGNED                (pipe_rx0_chanisaligned                     ),
    .PIPERX1CHANISALIGNED                (pipe_rx1_chanisaligned                     ),
    .PIPERX2CHANISALIGNED                (pipe_rx2_chanisaligned                     ),
    .PIPERX3CHANISALIGNED                (pipe_rx3_chanisaligned                     ),
    .PIPERX4CHANISALIGNED                (pipe_rx4_chanisaligned                     ),
    .PIPERX5CHANISALIGNED                (pipe_rx5_chanisaligned                     ),
    .PIPERX6CHANISALIGNED                (pipe_rx6_chanisaligned                     ),
    .PIPERX7CHANISALIGNED                (pipe_rx7_chanisaligned                     ),
    .PIPERX0STATUS                       (pipe_rx0_status                            ),
    .PIPERX1STATUS                       (pipe_rx1_status                            ),
    .PIPERX2STATUS                       (pipe_rx2_status                            ),
    .PIPERX3STATUS                       (pipe_rx3_status                            ),
    .PIPERX4STATUS                       (pipe_rx4_status                            ),
    .PIPERX5STATUS                       (pipe_rx5_status                            ),
    .PIPERX6STATUS                       (pipe_rx6_status                            ),
    .PIPERX7STATUS                       (pipe_rx7_status                            ),
    .PIPERX0PHYSTATUS                    (pipe_rx0_phy_status                        ),
    .PIPERX1PHYSTATUS                    (pipe_rx1_phy_status                        ),
    .PIPERX2PHYSTATUS                    (pipe_rx2_phy_status                        ),
    .PIPERX3PHYSTATUS                    (pipe_rx3_phy_status                        ),
    .PIPERX4PHYSTATUS                    (pipe_rx4_phy_status                        ),
    .PIPERX5PHYSTATUS                    (pipe_rx5_phy_status                        ),
    .PIPERX6PHYSTATUS                    (pipe_rx6_phy_status                        ),
    .PIPERX7PHYSTATUS                    (pipe_rx7_phy_status                        ),
    .PIPERX0ELECIDLE                     (pipe_rx0_elec_idle                         ),
    .PIPERX1ELECIDLE                     (pipe_rx1_elec_idle                         ),
    .PIPERX2ELECIDLE                     (pipe_rx2_elec_idle                         ),
    .PIPERX3ELECIDLE                     (pipe_rx3_elec_idle                         ),
    .PIPERX4ELECIDLE                     (pipe_rx4_elec_idle                         ),
    .PIPERX5ELECIDLE                     (pipe_rx5_elec_idle                         ),
    .PIPERX6ELECIDLE                     (pipe_rx6_elec_idle                         ),
    .PIPERX7ELECIDLE                     (pipe_rx7_elec_idle                         ),
    .PIPECLK                             (pipe_clk                                   ),
    .USERCLK                             (user_clk                                   ),
    .USERCLK2                            (user_clk2                                  ),
`ifdef VALIDATION
    .USERCLKPREBUF                       (user_clk_prebuf                            ),
    .USERCLKPREBUFEN                     (user_clk_prebuf_en                         ),
`endif
`ifdef B_TESTMODE
    .USERCLKPREBUF                       (user_clk_prebuf                            ),
    .USERCLKPREBUFEN                     (user_clk_prebuf_en                         ),
    .SCANMODEN                           (scanmode_n                                 ),
    .SCANENABLEN                         (scanenable_n                               ),
    .EDTCLK                              (edt_clk                                    ),
    .EDTUPDATE                           (edt_update                                 ),
    .EDTBYPASS                           (edt_bypass                                 ),
    .EDTCONFIGURATION                    (edt_configuration                          ),
    .EDTSINGLEBYPASSCHAIN                (edt_single_bypass_chain                    ),
    .EDTCHANNELSIN1                      (edt_channels_in1                           ),
    .EDTCHANNELSIN2                      (edt_channels_in2                           ),
    .EDTCHANNELSIN3                      (edt_channels_in3                           ),
    .EDTCHANNELSIN4                      (edt_channels_in4                           ),
    .EDTCHANNELSIN5                      (edt_channels_in5                           ),
    .EDTCHANNELSIN6                      (edt_channels_in6                           ),
    .EDTCHANNELSIN7                      (edt_channels_in7                           ),
    .EDTCHANNELSIN8                      (edt_channels_in8                           ),
    .PMVENABLEN                          (pmv_enable_n                               ),
    .PMVSELECT                           (pmv_select                                 ),
    .PMVDIVIDE                           (pmv_divide                                 ),
`endif
//`ifdef SECUREIP
//    .GSR                                 (gsr                                        ),
//`endif
    .SYSRSTN                             (sys_rst_n                                  ),
    .CMRSTN                              (cm_rst_n                                   ),
    .CMSTICKYRSTN                        (cm_sticky_rst_n                            ),
    .FUNCLVLRSTN                         (func_lvl_rst_n                             ),
    .TLRSTN                              (tl_rst_n                                   ),
    .DLRSTN                              (dl_rst_n                                   ),
    .PLRSTN                              (pl_rst_n                                   ),
    .PLTRANSMITHOTRST                    (pl_transmit_hot_rst                        ),
    // Global pins not on Holistic       model
    //.CFGRESET                          (cfg_reset                                  ),
    //.GWE                               (gwe                                        ),
    //.GRESTORE                          (grestore                                   ),
    //.GHIGHB                            (ghigh_b                                    ),
    .CFGMGMTDI                           (cfg_mgmt_di                                ),
    .CFGMGMTBYTEENN                      (cfg_mgmt_byte_en_n                         ),
    .CFGMGMTDWADDR                       (cfg_mgmt_dwaddr                            ),
    .CFGMGMTWRRW1CASRWN                  (cfg_mgmt_wr_rw1c_as_rw_n                   ),
    .CFGMGMTWRREADONLYN                  (cfg_mgmt_wr_readonly_n                     ),
    .CFGMGMTWRENN                        (cfg_mgmt_wr_en_n                           ),
    .CFGMGMTRDENN                        (cfg_mgmt_rd_en_n                           ),
    .CFGERRMALFORMEDN                    (cfg_err_malformed_n                        ),
    .CFGERRCORN                          (cfg_err_cor_n                              ),
    .CFGERRURN                           (cfg_err_ur_n                               ),
    .CFGERRECRCN                         (cfg_err_ecrc_n                             ),
    .CFGERRCPLTIMEOUTN                   (cfg_err_cpl_timeout_n                      ),
    .CFGERRCPLABORTN                     (cfg_err_cpl_abort_n                        ),
    .CFGERRCPLUNEXPECTN                  (cfg_err_cpl_unexpect_n                     ),
    .CFGERRPOISONEDN                     (cfg_err_poisoned_n                         ),
    .CFGERRACSN                          (cfg_err_acs_n                              ),
    .CFGERRATOMICEGRESSBLOCKEDN          (cfg_err_atomic_egress_blocked_n            ),
    .CFGERRMCBLOCKEDN                    (cfg_err_mc_blocked_n                       ),
    .CFGERRINTERNALUNCORN                (cfg_err_internal_uncor_n                   ),
    .CFGERRINTERNALCORN                  (cfg_err_internal_cor_n                     ),
    .CFGERRPOSTEDN                       (cfg_err_posted_n                           ),
    .CFGERRLOCKEDN                       (cfg_err_locked_n                           ),
    .CFGERRNORECOVERYN                   (cfg_err_norecovery_n                       ),
    .CFGERRAERHEADERLOG                  (cfg_err_aer_headerlog                      ),
    .CFGERRTLPCPLHEADER                  (cfg_err_tlp_cpl_header                     ),
    .CFGINTERRUPTN                       (cfg_interrupt_n                            ),
    .CFGINTERRUPTDI                      (cfg_interrupt_di                           ),
    .CFGINTERRUPTASSERTN                 (cfg_interrupt_assert_n                     ),
    .CFGINTERRUPTSTATN                   (cfg_interrupt_stat_n                       ),
    .CFGDSBUSNUMBER                      (cfg_ds_bus_number                          ),
    .CFGDSDEVICENUMBER                   (cfg_ds_device_number                       ),
    .CFGDSFUNCTIONNUMBER                 (cfg_ds_function_number                     ),
    .CFGPORTNUMBER                       (cfg_port_number                            ),
    .CFGPMHALTASPML0SN                   (cfg_pm_halt_aspm_l0s_n                     ),
    .CFGPMHALTASPML1N                    (cfg_pm_halt_aspm_l1_n                      ),
    .CFGPMFORCESTATEENN                  (cfg_pm_force_state_en_n                    ),
    .CFGPMFORCESTATE                     (cfg_pm_force_state                         ),
    .CFGPMWAKEN                          (cfg_pm_wake_n                              ),
    .CFGPMTURNOFFOKN                     (cfg_pm_turnoff_ok_n                        ),
    .CFGPMSENDPMETON                     (cfg_pm_send_pme_to_n                       ),
    .CFGPCIECAPINTERRUPTMSGNUM           (cfg_pciecap_interrupt_msgnum               ),
    .CFGTRNPENDINGN                      (cfg_trn_pending_n                          ),
    .CFGFORCEMPS                         (cfg_force_mps                              ),
    .CFGFORCECOMMONCLOCKOFF              (cfg_force_common_clock_off                 ),
    .CFGFORCEEXTENDEDSYNCON              (cfg_force_extended_sync_on                 ),
    .CFGDSN                              (cfg_dsn                                    ),
    .CFGDEVID                            (cfg_dev_id                                 ),
    .CFGVENDID                           (cfg_vend_id                                ),
    .CFGREVID                            (cfg_rev_id                                 ),
    .CFGSUBSYSID                         (cfg_subsys_id                              ),
    .CFGSUBSYSVENDID                     (cfg_subsys_vend_id                         ),
    .CFGAERINTERRUPTMSGNUM               (cfg_aer_interrupt_msgnum                   ),
    .DRPCLK                              (drp_clk                                    ),
    .DRPEN                               (drp_en                                     ),
    .DRPWE                               (drp_we                                     ),
    .DRPADDR                             (drp_addr                                   ),
    .DRPDI                               (drp_di                                     ),
    //.DRPREADPORT0                      (drp_read_port_0                            ),
    //.DRPREADPORT1                      (drp_read_port_1                            ),
    //.DRPREADPORT2                      (drp_read_port_2                            ),
    //.DRPREADPORT3                      (drp_read_port_3                            ),
    //.DRPREADPORT4                      (drp_read_port_4                            ),
    //.DRPREADPORT5                      (drp_read_port_5                            ),
    //.DRPREADPORT6                      (drp_read_port_6                            ),
    //.DRPREADPORT7                      (drp_read_port_7                            ),
    //.DRPREADPORT8                      (drp_read_port_8                            ),
    //.DRPREADPORT9                      (drp_read_port_9                            ),
    //.DRPREADPORT10                     (drp_read_port_10                           ),
    //.DRPREADPORT11                     (drp_read_port_11                           ),
    //.DRPREADPORT12                     (drp_read_port_12                           ),
    .DBGMODE                             (dbg_mode                                   ),
    .DBGSUBMODE                          (dbg_sub_mode                               ),
    .PLDBGMODE                           (pl_dbg_mode                                ),

    .TRNTDSTRDY                          (trn_tdst_rdy_bus                           ),
    .TRNTERRDROP                         (trn_terr_drop                              ),
    .TRNTBUFAV                           (trn_tbuf_av                                ),
    .TRNTCFGREQ                          (trn_tcfg_req                               ),
    .TRNRD                               (trn_rd                                     ),
    .TRNRREM                             (trn_rrem                                   ),
    .TRNRSOF                             (trn_rsof                                   ),
    .TRNREOF                             (trn_reof                                   ),
    .TRNRSRCRDY                          (trn_rsrc_rdy                               ),
    .TRNRSRCDSC                          (trn_rsrc_dsc                               ),
    .TRNRECRCERR                         (trn_recrc_err                              ),
    .TRNRERRFWD                          (trn_rerrfwd                                ),
    .TRNRBARHIT                          (trn_rbar_hit                               ),
    .TRNLNKUP                            (trn_lnk_up                                 ),
    .TRNFCPH                             (trn_fc_ph                                  ),
    .TRNFCPD                             (trn_fc_pd                                  ),
    .TRNFCNPH                            (trn_fc_nph                                 ),
    .TRNFCNPD                            (trn_fc_npd                                 ),
    .TRNFCCPLH                           (trn_fc_cplh                                ),
    .TRNFCCPLD                           (trn_fc_cpld                                ),
    .MIMTXWDATA                          (mim_tx_wdata                               ),
    .MIMTXWADDR                          (mim_tx_waddr                               ),
    .MIMTXWEN                            (mim_tx_wen                                 ),
    .MIMTXRADDR                          (mim_tx_raddr                               ),
    .MIMTXREN                            (mim_tx_ren                                 ),
    .MIMRXWDATA                          (mim_rx_wdata                               ),
    .MIMRXWADDR                          (mim_rx_waddr                               ),
    .MIMRXWEN                            (mim_rx_wen                                 ),
    .MIMRXRADDR                          (mim_rx_raddr                               ),
    .MIMRXREN                            (mim_rx_ren                                 ),
    .TRNTDLLPDSTRDY                      (trn_tdllp_dst_rdy                          ),
    .TRNRDLLPDATA                        (trn_rdllp_data                             ),
    .TRNRDLLPSRCRDY                      (trn_rdllp_src_rdy                          ),
    .LL2TFCINIT1SEQ                      (ll2_tfc_init1_seq                          ),
    .LL2TFCINIT2SEQ                      (ll2_tfc_init2_seq                          ),
    .PL2SUSPENDOK                        (pl2_suspend_ok                             ),
    .PL2RECOVERY                         (pl2_recovery                               ),
    .PL2RXELECIDLE                       (pl2_rx_elec_idle                           ),
    .PL2RXPMSTATE                        (pl2_rx_pm_state                            ),
    .PL2L0REQ                            (pl2_l0_req                                 ),
    .LL2SUSPENDOK                        (ll2_suspend_ok                             ),
    .LL2TXIDLE                           (ll2_tx_idle                                ),
    .LL2LINKSTATUS                       (ll2_link_status                            ),
    .TL2PPMSUSPENDOK                     (tl2_ppm_suspend_ok                         ),
    .TL2ASPMSUSPENDREQ                   (tl2_aspm_suspend_req                       ),
    .TL2ASPMSUSPENDCREDITCHECKOK         (tl2_aspm_suspend_credit_check_ok           ),
    .PL2LINKUP                           (pl2_link_up                                ),
    .PL2RECEIVERERR                      (pl2_receiver_err                           ),
    .LL2RECEIVERERR                      (ll2_receiver_err                           ),
    .LL2PROTOCOLERR                      (ll2_protocol_err                           ),
    .LL2BADTLPERR                        (ll2_bad_tlp_err                            ),
    .LL2BADDLLPERR                       (ll2_bad_dllp_err                           ),
    .LL2REPLAYROERR                      (ll2_replay_ro_err                          ),
    .LL2REPLAYTOERR                      (ll2_replay_to_err                          ),
    .TL2ERRHDR                           (tl2_err_hdr                                ),
    .TL2ERRMALFORMED                     (tl2_err_malformed                          ),
    .TL2ERRRXOVERFLOW                    (tl2_err_rxoverflow                         ),
    .TL2ERRFCPE                          (tl2_err_fcpe                               ),
    .PLSELLNKRATE                        (pl_sel_lnk_rate                            ),
    .PLSELLNKWIDTH                       (pl_sel_lnk_width                           ),
    .PLLTSSMSTATE                        (pl_ltssm_state                             ),
    .PLLANEREVERSALMODE                  (pl_lane_reversal_mode                      ),
    .PLPHYLNKUPN                         (pl_phy_lnk_up_n                            ),
    .PLTXPMSTATE                         (pl_tx_pm_state                             ),
    .PLRXPMSTATE                         (pl_rx_pm_state                             ),
    .PLLINKUPCFGCAP                      (pl_link_upcfg_cap                          ),
    .PLLINKGEN2CAP                       (pl_link_gen2_cap                           ),
    .PLLINKPARTNERGEN2SUPPORTED          (pl_link_partner_gen2_supported             ),
    .PLINITIALLINKWIDTH                  (pl_initial_link_width                      ),
    .PLDIRECTEDCHANGEDONE                (pl_directed_change_done                    ),
    .PIPETXRCVRDET                       (pipe_tx_rcvr_det                           ),
    .PIPETXRESET                         (pipe_tx_reset                              ),
    .PIPETXRATE                          (pipe_tx_rate                               ),
    .PIPETXDEEMPH                        (pipe_tx_deemph                             ),
    .PIPETXMARGIN                        (pipe_tx_margin                             ),
    .PIPERX0POLARITY                     (pipe_rx0_polarity                          ),
    .PIPERX1POLARITY                     (pipe_rx1_polarity                          ),
    .PIPERX2POLARITY                     (pipe_rx2_polarity                          ),
    .PIPERX3POLARITY                     (pipe_rx3_polarity                          ),
    .PIPERX4POLARITY                     (pipe_rx4_polarity                          ),
    .PIPERX5POLARITY                     (pipe_rx5_polarity                          ),
    .PIPERX6POLARITY                     (pipe_rx6_polarity                          ),
    .PIPERX7POLARITY                     (pipe_rx7_polarity                          ),
    .PIPETX0COMPLIANCE                   (pipe_tx0_compliance                        ),
    .PIPETX1COMPLIANCE                   (pipe_tx1_compliance                        ),
    .PIPETX2COMPLIANCE                   (pipe_tx2_compliance                        ),
    .PIPETX3COMPLIANCE                   (pipe_tx3_compliance                        ),
    .PIPETX4COMPLIANCE                   (pipe_tx4_compliance                        ),
    .PIPETX5COMPLIANCE                   (pipe_tx5_compliance                        ),
    .PIPETX6COMPLIANCE                   (pipe_tx6_compliance                        ),
    .PIPETX7COMPLIANCE                   (pipe_tx7_compliance                        ),
    .PIPETX0CHARISK                      (pipe_tx0_char_is_k                         ),
    .PIPETX1CHARISK                      (pipe_tx1_char_is_k                         ),
    .PIPETX2CHARISK                      (pipe_tx2_char_is_k                         ),
    .PIPETX3CHARISK                      (pipe_tx3_char_is_k                         ),
    .PIPETX4CHARISK                      (pipe_tx4_char_is_k                         ),
    .PIPETX5CHARISK                      (pipe_tx5_char_is_k                         ),
    .PIPETX6CHARISK                      (pipe_tx6_char_is_k                         ),
    .PIPETX7CHARISK                      (pipe_tx7_char_is_k                         ),
    .PIPETX0DATA                         (pipe_tx0_data                              ),
    .PIPETX1DATA                         (pipe_tx1_data                              ),
    .PIPETX2DATA                         (pipe_tx2_data                              ),
    .PIPETX3DATA                         (pipe_tx3_data                              ),
    .PIPETX4DATA                         (pipe_tx4_data                              ),
    .PIPETX5DATA                         (pipe_tx5_data                              ),
    .PIPETX6DATA                         (pipe_tx6_data                              ),
    .PIPETX7DATA                         (pipe_tx7_data                              ),
    .PIPETX0ELECIDLE                     (pipe_tx0_elec_idle                         ),
    .PIPETX1ELECIDLE                     (pipe_tx1_elec_idle                         ),
    .PIPETX2ELECIDLE                     (pipe_tx2_elec_idle                         ),
    .PIPETX3ELECIDLE                     (pipe_tx3_elec_idle                         ),
    .PIPETX4ELECIDLE                     (pipe_tx4_elec_idle                         ),
    .PIPETX5ELECIDLE                     (pipe_tx5_elec_idle                         ),
    .PIPETX6ELECIDLE                     (pipe_tx6_elec_idle                         ),
    .PIPETX7ELECIDLE                     (pipe_tx7_elec_idle                         ),
    .PIPETX0POWERDOWN                    (pipe_tx0_powerdown                         ),
    .PIPETX1POWERDOWN                    (pipe_tx1_powerdown                         ),
    .PIPETX2POWERDOWN                    (pipe_tx2_powerdown                         ),
    .PIPETX3POWERDOWN                    (pipe_tx3_powerdown                         ),
    .PIPETX4POWERDOWN                    (pipe_tx4_powerdown                         ),
    .PIPETX5POWERDOWN                    (pipe_tx5_powerdown                         ),
    .PIPETX6POWERDOWN                    (pipe_tx6_powerdown                         ),
    .PIPETX7POWERDOWN                    (pipe_tx7_powerdown                         ),
`ifdef B_TESTMODE
    .PMVOUT                              (pmv_out                                    ),
    .SCANOUT                             (scanout                                    ),
`endif
    .USERRSTN                            (user_rst_n                                 ),
    .PLRECEIVEDHOTRST                    (pl_received_hot_rst                        ),
    .RECEIVEDFUNCLVLRSTN                 (received_func_lvl_rst_n                    ),
    .LNKCLKEN                            (lnk_clk_en                                 ),
    .CFGMGMTDO                           (cfg_mgmt_do                                ),
    .CFGMGMTRDWRDONEN                    (cfg_mgmt_rd_wr_done_n                      ),
    .CFGERRAERHEADERLOGSETN              (cfg_err_aer_headerlog_set_n                ),
    .CFGERRCPLRDYN                       (cfg_err_cpl_rdy_n                          ),
    .CFGINTERRUPTRDYN                    (cfg_interrupt_rdy_n                        ),
    .CFGINTERRUPTMMENABLE                (cfg_interrupt_mmenable                     ),
    .CFGINTERRUPTMSIENABLE               (cfg_interrupt_msienable                    ),
    .CFGINTERRUPTDO                      (cfg_interrupt_do                           ),
    .CFGINTERRUPTMSIXENABLE              (cfg_interrupt_msixenable                   ),
    .CFGINTERRUPTMSIXFM                  (cfg_interrupt_msixfm                       ),
    .CFGMSGRECEIVED                      (cfg_msg_received                           ),
    .CFGMSGDATA                          (cfg_msg_data                               ),
    .CFGMSGRECEIVEDERRCOR                (cfg_msg_received_err_cor                   ),
    .CFGMSGRECEIVEDERRNONFATAL           (cfg_msg_received_err_non_fatal             ),
    .CFGMSGRECEIVEDERRFATAL              (cfg_msg_received_err_fatal                 ),
    .CFGMSGRECEIVEDASSERTINTA            (cfg_msg_received_assert_int_a              ),
    .CFGMSGRECEIVEDDEASSERTINTA          (cfg_msg_received_deassert_int_a            ),
    .CFGMSGRECEIVEDASSERTINTB            (cfg_msg_received_assert_int_b              ),
    .CFGMSGRECEIVEDDEASSERTINTB          (cfg_msg_received_deassert_int_b            ),
    .CFGMSGRECEIVEDASSERTINTC            (cfg_msg_received_assert_int_c              ),
    .CFGMSGRECEIVEDDEASSERTINTC          (cfg_msg_received_deassert_int_c            ),
    .CFGMSGRECEIVEDASSERTINTD            (cfg_msg_received_assert_int_d              ),
    .CFGMSGRECEIVEDDEASSERTINTD          (cfg_msg_received_deassert_int_d            ),
    .CFGMSGRECEIVEDPMPME                 (cfg_msg_received_pm_pme                    ),
    .CFGMSGRECEIVEDPMETOACK              (cfg_msg_received_pme_to_ack                ),
    .CFGMSGRECEIVEDPMETO                 (cfg_msg_received_pme_to                    ),
    .CFGMSGRECEIVEDSETSLOTPOWERLIMIT     (cfg_msg_received_setslotpowerlimit         ),
    .CFGMSGRECEIVEDUNLOCK                (cfg_msg_received_unlock                    ),
    .CFGMSGRECEIVEDPMASNAK               (cfg_msg_received_pm_as_nak                 ),
    .CFGPCIELINKSTATE                    (cfg_pcie_link_state                        ),
    .CFGPMRCVASREQL1N                    (cfg_pm_rcv_as_req_l1_n                     ),
    .CFGPMRCVREQACKN                     (cfg_pm_rcv_req_ack_n                       ),
    .CFGPMRCVENTERL1N                    (cfg_pm_rcv_enter_l1_n                      ),
    .CFGPMRCVENTERL23N                   (cfg_pm_rcv_enter_l23_n                     ),
    .CFGPMCSRPOWERSTATE                  (cfg_pmcsr_powerstate                       ),
    .CFGPMCSRPMEEN                       (cfg_pmcsr_pme_en                           ),
    .CFGPMCSRPMESTATUS                   (cfg_pmcsr_pme_status                       ),
    .CFGTRANSACTION                      (cfg_transaction                            ),
    .CFGTRANSACTIONTYPE                  (cfg_transaction_type                       ),
    .CFGTRANSACTIONADDR                  (cfg_transaction_addr                       ),
    .CFGCOMMANDIOENABLE                  (cfg_command_io_enable                      ),
    .CFGCOMMANDMEMENABLE                 (cfg_command_mem_enable                     ),
    .CFGCOMMANDBUSMASTERENABLE           (cfg_command_bus_master_enable              ),
    .CFGCOMMANDINTERRUPTDISABLE          (cfg_command_interrupt_disable              ),
    .CFGCOMMANDSERREN                    (cfg_command_serr_en                        ),
    .CFGBRIDGESERREN                     (cfg_bridge_serr_en                         ),
    .CFGDEVSTATUSCORRERRDETECTED         (cfg_dev_status_corr_err_detected           ),
    .CFGDEVSTATUSNONFATALERRDETECTED     (cfg_dev_status_non_fatal_err_detected      ),
    .CFGDEVSTATUSFATALERRDETECTED        (cfg_dev_status_fatal_err_detected          ),
    .CFGDEVSTATUSURDETECTED              (cfg_dev_status_ur_detected                 ),
    .CFGDEVCONTROLCORRERRREPORTINGEN     (cfg_dev_control_corr_err_reporting_en      ),
    .CFGDEVCONTROLNONFATALREPORTINGEN    (cfg_dev_control_non_fatal_reporting_en     ),
    .CFGDEVCONTROLFATALERRREPORTINGEN    (cfg_dev_control_fatal_err_reporting_en     ),
    .CFGDEVCONTROLURERRREPORTINGEN       (cfg_dev_control_ur_err_reporting_en        ),
    .CFGDEVCONTROLENABLERO               (cfg_dev_control_enable_ro                  ),
    .CFGDEVCONTROLMAXPAYLOAD             (cfg_dev_control_max_payload                ),
    .CFGDEVCONTROLEXTTAGEN               (cfg_dev_control_ext_tag_en                 ),
    .CFGDEVCONTROLPHANTOMEN              (cfg_dev_control_phantom_en                 ),
    .CFGDEVCONTROLAUXPOWEREN             (cfg_dev_control_aux_power_en               ),
    .CFGDEVCONTROLNOSNOOPEN              (cfg_dev_control_no_snoop_en                ),
    .CFGDEVCONTROLMAXREADREQ             (cfg_dev_control_max_read_req               ),
    .CFGLINKSTATUSCURRENTSPEED           (cfg_link_status_current_speed              ),
    .CFGLINKSTATUSNEGOTIATEDWIDTH        (cfg_link_status_negotiated_width           ),
    .CFGLINKSTATUSLINKTRAINING           (cfg_link_status_link_training              ),
    .CFGLINKSTATUSDLLACTIVE              (cfg_link_status_dll_active                 ),
    .CFGLINKSTATUSBANDWIDTHSTATUS        (cfg_link_status_bandwidth_status           ),
    .CFGLINKSTATUSAUTOBANDWIDTHSTATUS    (cfg_link_status_auto_bandwidth_status      ),
    .CFGLINKCONTROLASPMCONTROL           (cfg_link_control_aspm_control              ),
    .CFGLINKCONTROLRCB                   (cfg_link_control_rcb                       ),
    .CFGLINKCONTROLLINKDISABLE           (cfg_link_control_link_disable              ),
    .CFGLINKCONTROLRETRAINLINK           (cfg_link_control_retrain_link              ),
    .CFGLINKCONTROLCOMMONCLOCK           (cfg_link_control_common_clock              ),
    .CFGLINKCONTROLEXTENDEDSYNC          (cfg_link_control_extended_sync             ),
    .CFGLINKCONTROLCLOCKPMEN             (cfg_link_control_clock_pm_en               ),
    .CFGLINKCONTROLHWAUTOWIDTHDIS        (cfg_link_control_hw_auto_width_dis         ),
    .CFGLINKCONTROLBANDWIDTHINTEN        (cfg_link_control_bandwidth_int_en          ),
    .CFGLINKCONTROLAUTOBANDWIDTHINTEN    (cfg_link_control_auto_bandwidth_int_en     ),
    .CFGDEVCONTROL2CPLTIMEOUTVAL         (cfg_dev_control2_cpl_timeout_val           ),
    .CFGDEVCONTROL2CPLTIMEOUTDIS         (cfg_dev_control2_cpl_timeout_dis           ),
    .CFGDEVCONTROL2ARIFORWARDEN          (cfg_dev_control2_ari_forward_en            ),
    .CFGDEVCONTROL2ATOMICREQUESTEREN     (cfg_dev_control2_atomic_requester_en       ),
    .CFGDEVCONTROL2ATOMICEGRESSBLOCK     (cfg_dev_control2_atomic_egress_block       ),
    .CFGDEVCONTROL2IDOREQEN              (cfg_dev_control2_ido_req_en                ),
    .CFGDEVCONTROL2IDOCPLEN              (cfg_dev_control2_ido_cpl_en                ),
    .CFGDEVCONTROL2LTREN                 (cfg_dev_control2_ltr_en                    ),
    .CFGDEVCONTROL2TLPPREFIXBLOCK        (cfg_dev_control2_tlp_prefix_block          ),
    .CFGSLOTCONTROLELECTROMECHILCTLPULSE (cfg_slot_control_electromech_il_ctl_pulse  ),
    .CFGROOTCONTROLSYSERRCORRERREN       (cfg_root_control_syserr_corr_err_en        ),
    .CFGROOTCONTROLSYSERRNONFATALERREN   (cfg_root_control_syserr_non_fatal_err_en   ),
    .CFGROOTCONTROLSYSERRFATALERREN      (cfg_root_control_syserr_fatal_err_en       ),
    .CFGROOTCONTROLPMEINTEN              (cfg_root_control_pme_int_en                ),
    .CFGAERECRCCHECKEN                   (cfg_aer_ecrc_check_en                      ),
    .CFGAERECRCGENEN                     (cfg_aer_ecrc_gen_en                        ),
    .CFGAERROOTERRCORRERRREPORTINGEN     (cfg_aer_rooterr_corr_err_reporting_en      ),
    .CFGAERROOTERRNONFATALERRREPORTINGEN (cfg_aer_rooterr_non_fatal_err_reporting_en ),
    .CFGAERROOTERRFATALERRREPORTINGEN    (cfg_aer_rooterr_fatal_err_reporting_en     ),
    .CFGAERROOTERRCORRERRRECEIVED        (cfg_aer_rooterr_corr_err_received          ),
    .CFGAERROOTERRNONFATALERRRECEIVED    (cfg_aer_rooterr_non_fatal_err_received     ),
    .CFGAERROOTERRFATALERRRECEIVED       (cfg_aer_rooterr_fatal_err_received         ),
    .CFGVCTCVCMAP                        (cfg_vc_tcvc_map                            ),
    .DRPRDY                              (drp_rdy                                    ),
    .DRPDO                               (drp_do                                     ),
    //.DRPWRITEEN                        (drp_write_en                               ),
    //.DRPWRITEPORT0                     (drp_write_port_0                           ),
    //.DRPWRITEPORT1                     (drp_write_port_1                           ),
    //.DRPWRITEPORT2                     (drp_write_port_2                           ),
    //.DRPWRITEPORT3                     (drp_write_port_3                           ),
    //.DRPWRITEPORT4                     (drp_write_port_4                           ),
    //.DRPWRITEPORT5                     (drp_write_port_5                           ),
    //.DRPWRITEPORT6                     (drp_write_port_6                           ),
    //.DRPWRITEPORT7                     (drp_write_port_7                           ),
    //.DRPWRITEPORT8                     (drp_write_port_8                           ),
    //.DRPWRITEPORT9                     (drp_write_port_9                           ),
    //.DRPWRITEPORT10                    (drp_write_port_10                          ),
    //.DRPWRITEPORT11                    (drp_write_port_11                          ),
    //.DRPWRITEPORT12                    (drp_write_port_12                          ),
    //.DRPREADADDR                       (drp_read_addr                              ),
    .DBGVECA                             (dbg_vec_a                                  ),
    .DBGVECB                             (dbg_vec_b                                  ),
    .DBGVECC                             (dbg_vec_c                                  ),
    .DBGSCLRA                            (dbg_sclr_a                                 ),
    .DBGSCLRB                            (dbg_sclr_b                                 ),
    .DBGSCLRC                            (dbg_sclr_c                                 ),
    .DBGSCLRD                            (dbg_sclr_d                                 ),
    .DBGSCLRE                            (dbg_sclr_e                                 ),
    .DBGSCLRF                            (dbg_sclr_f                                 ),
    .DBGSCLRG                            (dbg_sclr_g                                 ),
    .DBGSCLRH                            (dbg_sclr_h                                 ),
    .DBGSCLRI                            (dbg_sclr_i                                 ),
    .DBGSCLRJ                            (dbg_sclr_j                                 ),
    .DBGSCLRK                            (dbg_sclr_k                                 ),
    .PLDBGVEC                            (pl_dbg_vec                                 )
    //.XILUNCONNOUT                      (xil_unconn_out                             )
  );
endmodule




`timescale 1ns/1ps
module model_ap2_tst_pcie_bram_top_7x
#(
  parameter IMPL_TARGET               = "HARD",        // the implementation target : HARD, SOFT
  parameter DEV_CAP_MAX_PAYLOAD_SUPPORTED = 0,         // MPS Supported : 0 - 128 B, 1 - 256 B, 2 - 512 B, 3 - 1024 B
  parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,     // PCIe Link Speed : 1 - 2.5 GT/s; 2 - 5.0 GT/s
  parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,    // PCIe Link Width : 1 / 2 / 4 / 8

  parameter VC0_TX_LASTPACKET         = 31,            // Number of Packets in Transmit
  parameter TLM_TX_OVERHEAD           = 24,            // Overhead Bytes for Packets (Transmit)
  parameter TL_TX_RAM_RADDR_LATENCY   = 1,             // BRAM Read Address Latency (Transmit)
  parameter TL_TX_RAM_RDATA_LATENCY   = 2,             // BRAM Read Data Latency (Transmit)
  parameter TL_TX_RAM_WRITE_LATENCY   = 1,             // BRAM Write Latency (Transmit)

  parameter VC0_RX_RAM_LIMIT          = 'h1FFF,        // RAM Size (Receive)
  parameter TL_RX_RAM_RADDR_LATENCY   = 1,             // BRAM Read Address Latency (Receive)
  parameter TL_RX_RAM_RDATA_LATENCY   = 2,             // BRAM Read Data Latency (Receive)
  parameter TL_RX_RAM_WRITE_LATENCY   = 1              // BRAM Write Latency (Receive)
)
(
  input          user_clk_i,                  // Clock input
  input          reset_i,                     // Reset input

  input          mim_tx_wen,                  // Write Enable for Transmit path BRAM
  input  [12:0]  mim_tx_waddr,                // Write Address for Transmit path BRAM
  input  [71:0]  mim_tx_wdata,                // Write Data for Transmit path BRAM
  input          mim_tx_ren,                  // Read Enable for Transmit path BRAM
  input          mim_tx_rce,                  // Read Output Register Clock Enable for Transmit path BRAM
  input  [12:0]  mim_tx_raddr,                // Read Address for Transmit path BRAM
  output [71:0]  mim_tx_rdata,                // Read Data for Transmit path BRAM

  input          mim_rx_wen,                  // Write Enable for Receive path BRAM
  input  [12:0]  mim_rx_waddr,                // Write Enable for Receive path BRAM
  input  [71:0]  mim_rx_wdata,                // Write Enable for Receive path BRAM
  input          mim_rx_ren,                  // Read Enable for Receive path BRAM
  input          mim_rx_rce,                  // Read Output Register Clock Enable for Receive path BRAM
  input  [12:0]  mim_rx_raddr,                // Read Address for Receive path BRAM
  output [71:0]  mim_rx_rdata                 // Read Data for Receive path BRAM
);

  // TX calculations
  localparam MPS_BYTES = ((DEV_CAP_MAX_PAYLOAD_SUPPORTED == 0) ? 128 :
                          (DEV_CAP_MAX_PAYLOAD_SUPPORTED == 1) ? 256 :
                          (DEV_CAP_MAX_PAYLOAD_SUPPORTED == 2) ? 512 :
                                                                1024 );

  localparam BYTES_TX = (VC0_TX_LASTPACKET + 1) * (MPS_BYTES + TLM_TX_OVERHEAD);

  localparam ROWS_TX = 1;
  localparam COLS_TX = ((BYTES_TX <= 4096) ?  1 :
                        (BYTES_TX <= 8192) ?  2 :
                        (BYTES_TX <= 16384) ? 4 :
                        (BYTES_TX <= 32768) ? 8 :
                                             18
                       );

  // RX calculations
  localparam ROWS_RX = 1;

  localparam COLS_RX = ((VC0_RX_RAM_LIMIT < 'h0200) ? 1 :
                        (VC0_RX_RAM_LIMIT < 'h0400) ? 2 :
                        (VC0_RX_RAM_LIMIT < 'h0800) ? 4 :
                        (VC0_RX_RAM_LIMIT < 'h1000) ? 8 :
                                                 18
                       );

  initial begin
     $display("[%t] %m ROWS_TX %0d COLS_TX %0d", $time, ROWS_TX, COLS_TX);
     $display("[%t] %m ROWS_RX %0d COLS_RX %0d", $time, ROWS_RX, COLS_RX);
  end

model_ap2_tst_pcie_brams_7x #(
    .LINK_CAP_MAX_LINK_WIDTH ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_MAX_LINK_SPEED ( LINK_CAP_MAX_LINK_SPEED ),
    .IMPL_TARGET             ( IMPL_TARGET ),
    .NUM_BRAMS               ( COLS_TX ),
    .RAM_RADDR_LATENCY       ( TL_TX_RAM_RADDR_LATENCY ),
    .RAM_RDATA_LATENCY       ( TL_TX_RAM_RDATA_LATENCY ),
    .RAM_WRITE_LATENCY       ( TL_TX_RAM_WRITE_LATENCY )
  ) 
  model_ap2_tst_pcie_brams_tx (
    .user_clk_i ( user_clk_i ),
    .reset_i    ( reset_i ),
    .waddr      ( mim_tx_waddr ),
    .wen        ( mim_tx_wen ),
    .ren        ( mim_tx_ren ),
    .rce        ( mim_tx_rce ),
    .wdata      ( mim_tx_wdata ),
    .raddr      ( mim_tx_raddr ),
    .rdata      ( mim_tx_rdata )
  );

model_ap2_tst_pcie_brams_7x #(
    .LINK_CAP_MAX_LINK_WIDTH ( LINK_CAP_MAX_LINK_WIDTH ),
    .LINK_CAP_MAX_LINK_SPEED ( LINK_CAP_MAX_LINK_SPEED ),
    .IMPL_TARGET             ( IMPL_TARGET ),
    .NUM_BRAMS               ( COLS_RX ),
    .RAM_RADDR_LATENCY       ( TL_RX_RAM_RADDR_LATENCY ),
    .RAM_RDATA_LATENCY       ( TL_RX_RAM_RDATA_LATENCY ),
    .RAM_WRITE_LATENCY       ( TL_RX_RAM_WRITE_LATENCY )
  ) model_ap2_tst_pcie_brams_rx (
    .user_clk_i ( user_clk_i ),
    .reset_i    ( reset_i ),
    .waddr      ( mim_rx_waddr ),
    .wen        ( mim_rx_wen ),
    .ren        ( mim_rx_ren ),
    .rce        ( mim_rx_rce ),
    .wdata      ( mim_rx_wdata ),
    .raddr      ( mim_rx_raddr ),
    .rdata      ( mim_rx_rdata )
   );

endmodule // pcie_bram_top


`timescale 1ns/1ps
module model_ap2_tst_pcie_brams_7x
#(
  parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,        // PCIe Link Speed : 1 - 2.5 GT/s; 2 - 5.0 GT/s
  parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,       // PCIe Link Width : 1 / 2 / 4 / 8
  parameter IMPL_TARGET             = "HARD",             // the implementation target : HARD, SOFT

  // the number of BRAMs to use
  // supported values are:
  // 1,2,4,8,18
  parameter NUM_BRAMS               = 0,

  // BRAM read address latency
  //
  // value     meaning
  // ====================================================
  //   0       BRAM read address port sample
  //   1       BRAM read address port sample and a pipeline stage on the address port
  parameter RAM_RADDR_LATENCY   = 1,

  // BRAM read data latency
  //
  // value     meaning
  // ====================================================
  //   1       no BRAM OREG
  //   2       use BRAM OREG
  //   3       use BRAM OREG and a pipeline stage on the data port
  parameter RAM_RDATA_LATENCY   = 1,

  // BRAM write latency
  // The BRAM write port is synchronous
  //
  // value     meaning
  // ====================================================
  //   0       BRAM write port sample
  //   1       BRAM write port sample plus pipeline stage
  parameter RAM_WRITE_LATENCY       = 1,
  parameter TCQ           = 1 // synthesis warning removed: parameter declaration becomes local
)
(
  input          user_clk_i,
  input          reset_i,

  input          wen,
  input  [12:0]  waddr,
  input  [71:0]  wdata,
  input          ren,
  input          rce,
  input  [12:0]  raddr,
  output [71:0]  rdata
  );

  // turn on the bram output register
  localparam DOB_REG = (RAM_RDATA_LATENCY > 1) ? 1 : 0;

  // calculate the data width of the individual brams
  localparam [6:0] WIDTH = ((NUM_BRAMS == 1) ? 72 :
                            (NUM_BRAMS == 2) ? 36 :
                            (NUM_BRAMS == 4) ? 18 :
                            (NUM_BRAMS == 8) ?  9 :
                                                4
                           );

//  parameter TCQ           = 1;

  wire        wen_int;
  wire [12:0] waddr_int;
  wire [71:0] wdata_int;

  wire        ren_int;
  wire [12:0] raddr_int;
  wire [71:0] rdata_int;

  //synthesis translate_off
  initial
  begin
    $display("[%t] %m NUM_BRAMS %0d  DOB_REG %0d WIDTH %0d RAM_WRITE_LATENCY %0d RAM_RADDR_LATENCY %0d RAM_RDATA_LATENCY %0d",
    $time, NUM_BRAMS, DOB_REG, WIDTH, RAM_WRITE_LATENCY, RAM_RADDR_LATENCY, RAM_RDATA_LATENCY);

    case (NUM_BRAMS)
      1,2,4,8,18:;
      default:
        begin
           $display("[%t] %m Error NUM_BRAMS %0d not supported", $time, NUM_BRAMS);
           $finish;
        end
    endcase // case(NUM_BRAMS)

    case (RAM_RADDR_LATENCY)
      0,1:;
      default:
        begin
           $display("[%t] %m Error RAM_READ_LATENCY %0d not supported", $time, RAM_RADDR_LATENCY);
           $finish;
        end
    endcase // case (RAM_RADDR_LATENCY)

    case (RAM_RDATA_LATENCY)
      1,2,3:;
      default:
        begin
           $display("[%t] %m Error RAM_READ_LATENCY %0d not supported", $time, RAM_RDATA_LATENCY);
           $finish;
        end
    endcase // case (RAM_RDATA_LATENCY)

    case (RAM_WRITE_LATENCY)
      0,1:;
      default:
        begin
           $display("[%t] %m Error RAM_WRITE_LATENCY %0d not supported", $time, RAM_WRITE_LATENCY);
           $finish;
        end
    endcase // case(RAM_WRITE_LATENCY)

  end
  //synthesis translate_on

  // model the delays for ram write latency

  generate if (RAM_WRITE_LATENCY == 1) begin : wr_lat_2
   reg        wen_q;
   reg [12:0] waddr_q;
   reg [71:0] wdata_q;

    always @(posedge user_clk_i) begin
      if (reset_i)
      begin
        wen_q   <= #TCQ 1'b0;
        waddr_q <= #TCQ 13'b0;
      // Disable Reset on Data Path @ BRAM i/f as I/O come from PCIe HB.
      //  wdata_q <= #TCQ 72'b0;
      end 
      else 
      begin
        wen_q   <= #TCQ wen;
        waddr_q <= #TCQ waddr;
        wdata_q <= #TCQ wdata;
      end
    end

    assign wen_int   = wen_q;
    assign waddr_int = waddr_q;
    assign wdata_int = wdata_q;
  end // if (RAM_WRITE_LATENCY == 1)

  else if (RAM_WRITE_LATENCY == 0) begin : wr_lat_1
    assign wen_int   = wen;
    assign waddr_int = waddr;
    assign wdata_int = wdata;
  end
  endgenerate

  // model the delays for ram read latency

  generate if (RAM_RADDR_LATENCY == 1) begin : raddr_lat_2
    reg        ren_q;
    reg [12:0] raddr_q;

    always @(posedge user_clk_i) begin
      if (reset_i)
      begin
        ren_q   <= #TCQ 1'b0;
        raddr_q <= #TCQ 13'b0;
      end
      else
      begin
        ren_q   <= #TCQ ren;
        raddr_q <= #TCQ raddr;
      end // else: !if(reset_i)
    end

    assign ren_int   = ren_q;
    assign raddr_int = raddr_q;
  end // block: rd_lat_addr_2

  else begin : raddr_lat_1
    assign ren_int   = ren;
    assign raddr_int = raddr;
  end
  endgenerate

  generate if (RAM_RDATA_LATENCY == 3) begin : rdata_lat_3
    reg [71:0] rdata_q;

    always @(posedge user_clk_i) begin
      // Disable Reset on Data Path @ BRAM i/f as I/O come from PCIe HB.
      //if (reset_i)
      //begin
      //  rdata_q <= #TCQ 72'b0;
      //end
      //else
      //begin
        rdata_q <= #TCQ rdata_int;
      //end // else: !if(reset_i)
    end

    assign rdata     = rdata_q;

  end // block: rd_lat_data_3

  else begin : rdata_lat_1_2
    assign rdata     = rdata_int;
  end
  endgenerate

  // instantiate the brams
  generate
    genvar ii;
    for (ii = 0; ii < NUM_BRAMS; ii = ii + 1) begin : brams
model_ap2_tst_pcie_bram_7x #(
        .LINK_CAP_MAX_LINK_WIDTH(LINK_CAP_MAX_LINK_WIDTH),
        .LINK_CAP_MAX_LINK_SPEED(LINK_CAP_MAX_LINK_SPEED),
        .IMPL_TARGET      (IMPL_TARGET),
        .DOB_REG          (DOB_REG),
        .WIDTH            (WIDTH)
      )
      model_ap2_tst_ram (
        .user_clk_i(user_clk_i),
        .reset_i(reset_i),
        .wen_i(wen_int),
        .waddr_i(waddr_int),
        .wdata_i(wdata_int[(((ii + 1) * WIDTH) - 1): (ii * WIDTH)]),
        .ren_i(ren_int),
        .raddr_i(raddr_int),
        .rdata_o(rdata_int[(((ii + 1) * WIDTH) - 1): (ii * WIDTH)]),
        .rce_i(rce)
      );
    end
  endgenerate

endmodule // pcie_brams_7x



`timescale 1ns/1ps
module model_ap2_tst_pcie_bram_7x
  #(
    parameter [3:0]  LINK_CAP_MAX_LINK_SPEED = 4'h1,        // PCIe Link Speed : 1 - 2.5 GT/s; 2 - 5.0 GT/s
    parameter [5:0]  LINK_CAP_MAX_LINK_WIDTH = 6'h08,       // PCIe Link Width : 1 / 2 / 4 / 8
    parameter IMPL_TARGET = "HARD",                         // the implementation target : HARD, SOFT
    parameter DOB_REG = 0,                                  // 1 - use the output register;
                                                            // 0 - don't use the output register
    parameter WIDTH = 0                                     // supported WIDTH's : 4, 9, 18, 36 - uses RAMB36
                                                            //                     72 - uses RAMB36SDP
    )
    (
     input               user_clk_i,// user clock
     input               reset_i,   // bram reset

     input               wen_i,     // write enable
     input [12:0]        waddr_i,   // write address
     input [WIDTH - 1:0] wdata_i,   // write data

     input               ren_i,     // read enable
     input               rce_i,     // output register clock enable
     input [12:0]        raddr_i,   // read address

     output [WIDTH - 1:0] rdata_o   // read data
     );

   // map the address bits
   localparam ADDR_MSB = ((WIDTH == 4)  ? 12 :
                          (WIDTH == 9)  ? 11 :
                          (WIDTH == 18) ? 10 :
                          (WIDTH == 36) ?  9 :
                                           8
                          );

   // set the width of the tied off low address bits
   localparam ADDR_LO_BITS = ((WIDTH == 4)  ? 2 :
                              (WIDTH == 9)  ? 3 :
                              (WIDTH == 18) ? 4 :
                              (WIDTH == 36) ? 5 :
                                              0 // for WIDTH 72 use RAMB36SDP
                              );

   // map the data bits
   localparam D_MSB =  ((WIDTH == 4)  ?  3 :
                        (WIDTH == 9)  ?  7 :
                        (WIDTH == 18) ? 15 :
                        (WIDTH == 36) ? 31 :
                                        63
                        );

   // map the data parity bits
   localparam DP_LSB =  D_MSB + 1;

   localparam DP_MSB =  ((WIDTH == 4)  ? 4 :
                         (WIDTH == 9)  ? 8 :
                         (WIDTH == 18) ? 17 :
                         (WIDTH == 36) ? 35 :
                                         71
                        );

   localparam DPW = DP_MSB - DP_LSB + 1;
   localparam WRITE_MODE = ((WIDTH == 72) && (!((LINK_CAP_MAX_LINK_SPEED == 4'h2) && (LINK_CAP_MAX_LINK_WIDTH == 6'h08)))) ? "WRITE_FIRST" :
                           ((LINK_CAP_MAX_LINK_SPEED == 4'h2) && (LINK_CAP_MAX_LINK_WIDTH == 6'h08)) ? "WRITE_FIRST" : "NO_CHANGE";

   localparam DEVICE = (IMPL_TARGET == "HARD") ? "7SERIES" : "VIRTEX6";
   localparam BRAM_SIZE = "36Kb";

   localparam WE_WIDTH =(DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES") ?
                            ((WIDTH <= 9) ? 1 :
                             (WIDTH > 9 && WIDTH <= 18) ? 2 :
                             (WIDTH > 18 && WIDTH <= 36) ? 4 :
                             (WIDTH > 36 && WIDTH <= 72) ? 8 :
                             (BRAM_SIZE == "18Kb") ? 4 : 8 ) : 8;

   //synthesis translate_off
   initial begin
      //$display("[%t] %m DOB_REG %0d WIDTH %0d ADDR_MSB %0d ADDR_LO_BITS %0d DP_MSB %0d DP_LSB %0d D_MSB %0d",
      //          $time, DOB_REG,   WIDTH,    ADDR_MSB,    ADDR_LO_BITS,    DP_MSB,    DP_LSB,    D_MSB);

      case (WIDTH)
        4,9,18,36,72:;
        default:
          begin
             $display("[%t] %m Error WIDTH %0d not supported", $time, WIDTH);
             $finish;
          end
      endcase // case (WIDTH)
   end
   //synthesis translate_on

   generate
   if ((LINK_CAP_MAX_LINK_WIDTH == 6'h08 && LINK_CAP_MAX_LINK_SPEED == 4'h2) || (WIDTH == 72)) begin : use_sdp
        BRAM_SDP_MACRO_model #(
               .DEVICE        (DEVICE),
               .BRAM_SIZE     (BRAM_SIZE),
               .DO_REG        (DOB_REG),
               .READ_WIDTH    (WIDTH),
               .WRITE_WIDTH   (WIDTH),
               .WRITE_MODE    (WRITE_MODE)
               )
        ramb36sdp(
               .DO             (rdata_o[WIDTH-1:0]),
               .DI             (wdata_i[WIDTH-1:0]),
               .RDADDR         (raddr_i[ADDR_MSB:0]),
               .RDCLK          (user_clk_i),
               .RDEN           (ren_i),
               .REGCE          (rce_i),
               .RST            (reset_i),
               .WE             ({WE_WIDTH{1'b1}}),
               .WRADDR         (waddr_i[ADDR_MSB:0]),
               .WRCLK          (user_clk_i),
               .WREN           (wen_i)
               );

    end  // block: use_sdp
    else if (WIDTH <= 36) begin : use_tdp
    // use RAMB36's if the width is 4, 9, 18, or 36
        BRAM_TDP_MACRO #(
               .DEVICE        (DEVICE),
               .BRAM_SIZE     (BRAM_SIZE),
               .DOA_REG       (0),
               .DOB_REG       (DOB_REG),
               .READ_WIDTH_A  (WIDTH),
               .READ_WIDTH_B  (WIDTH),
               .WRITE_WIDTH_A (WIDTH),
               .WRITE_WIDTH_B (WIDTH),
               .WRITE_MODE_A  (WRITE_MODE)
               )
        ramb36(
               .DOA            (),
               .DOB            (rdata_o[WIDTH-1:0]),
               .ADDRA          (waddr_i[ADDR_MSB:0]),
               .ADDRB          (raddr_i[ADDR_MSB:0]),
               .CLKA           (user_clk_i),
               .CLKB           (user_clk_i),
               .DIA            (wdata_i[WIDTH-1:0]),
               .DIB            ({WIDTH{1'b0}}),
               .ENA            (wen_i),
               .ENB            (ren_i),
               .REGCEA         (1'b0),
               .REGCEB         (rce_i),
               .RSTA           (reset_i),
               .RSTB           (reset_i),
               .WEA            ({WE_WIDTH{1'b1}}),
               .WEB            ({WE_WIDTH{1'b0}})
               );
   end // block: use_tdp
   endgenerate

endmodule // pcie_bram_7x



`timescale 1ns/1ps
module model_ap2_tst_pcie_pipe_pipeline #
(
  parameter        LINK_CAP_MAX_LINK_WIDTH = 8,
  parameter        PIPE_PIPELINE_STAGES = 0    // 0 - 0 stages, 1 - 1 stage, 2 - 2 stages
)
(
  // Pipe Per-Link Signals
  input   wire        pipe_tx_rcvr_det_i       ,
  input   wire        pipe_tx_reset_i          ,
  input   wire        pipe_tx_rate_i           ,
  input   wire        pipe_tx_deemph_i         ,
  input   wire [2:0]  pipe_tx_margin_i         ,
  input   wire        pipe_tx_swing_i          ,

  output  wire        pipe_tx_rcvr_det_o       ,
  output  wire        pipe_tx_reset_o          ,
  output  wire        pipe_tx_rate_o           ,
  output  wire        pipe_tx_deemph_o         ,
  output  wire [2:0]  pipe_tx_margin_o         ,
  output  wire        pipe_tx_swing_o          ,

  // Pipe Per-Lane Signals - Lane 0
  output  wire [ 1:0] pipe_rx0_char_is_k_o     ,
  output  wire [15:0] pipe_rx0_data_o          ,
  output  wire        pipe_rx0_valid_o         ,
  output  wire        pipe_rx0_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx0_status_o        ,
  output  wire        pipe_rx0_phy_status_o    ,
  output  wire        pipe_rx0_elec_idle_o     ,
  input   wire        pipe_rx0_polarity_i      ,
  input   wire        pipe_tx0_compliance_i    ,
  input   wire [ 1:0] pipe_tx0_char_is_k_i     ,
  input   wire [15:0] pipe_tx0_data_i          ,
  input   wire        pipe_tx0_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx0_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx0_char_is_k_i     ,
  input  wire [15:0]  pipe_rx0_data_i         ,
  input  wire         pipe_rx0_valid_i         ,
  input  wire         pipe_rx0_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx0_status_i        ,
  input  wire         pipe_rx0_phy_status_i    ,
  input  wire         pipe_rx0_elec_idle_i     ,
  output wire         pipe_rx0_polarity_o      ,
  output wire         pipe_tx0_compliance_o    ,
  output wire [ 1:0]  pipe_tx0_char_is_k_o     ,
  output wire [15:0]  pipe_tx0_data_o          ,
  output wire         pipe_tx0_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx0_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 1
  output  wire [ 1:0] pipe_rx1_char_is_k_o     ,
  output  wire [15:0] pipe_rx1_data_o         ,
  output  wire        pipe_rx1_valid_o         ,
  output  wire        pipe_rx1_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx1_status_o        ,
  output  wire        pipe_rx1_phy_status_o    ,
  output  wire        pipe_rx1_elec_idle_o     ,
  input   wire        pipe_rx1_polarity_i      ,
  input   wire        pipe_tx1_compliance_i    ,
  input   wire [ 1:0] pipe_tx1_char_is_k_i     ,
  input   wire [15:0] pipe_tx1_data_i          ,
  input   wire        pipe_tx1_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx1_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx1_char_is_k_i     ,
  input  wire [15:0]  pipe_rx1_data_i         ,
  input  wire         pipe_rx1_valid_i         ,
  input  wire         pipe_rx1_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx1_status_i        ,
  input  wire         pipe_rx1_phy_status_i    ,
  input  wire         pipe_rx1_elec_idle_i     ,
  output wire         pipe_rx1_polarity_o      ,
  output wire         pipe_tx1_compliance_o    ,
  output wire [ 1:0]  pipe_tx1_char_is_k_o     ,
  output wire [15:0]  pipe_tx1_data_o          ,
  output wire         pipe_tx1_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx1_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 2
  output  wire [ 1:0] pipe_rx2_char_is_k_o     ,
  output  wire [15:0] pipe_rx2_data_o         ,
  output  wire        pipe_rx2_valid_o         ,
  output  wire        pipe_rx2_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx2_status_o        ,
  output  wire        pipe_rx2_phy_status_o    ,
  output  wire        pipe_rx2_elec_idle_o     ,
  input   wire        pipe_rx2_polarity_i      ,
  input   wire        pipe_tx2_compliance_i    ,
  input   wire [ 1:0] pipe_tx2_char_is_k_i     ,
  input   wire [15:0] pipe_tx2_data_i          ,
  input   wire        pipe_tx2_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx2_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx2_char_is_k_i     ,
  input  wire [15:0]  pipe_rx2_data_i         ,
  input  wire         pipe_rx2_valid_i         ,
  input  wire         pipe_rx2_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx2_status_i        ,
  input  wire         pipe_rx2_phy_status_i    ,
  input  wire         pipe_rx2_elec_idle_i     ,
  output wire         pipe_rx2_polarity_o      ,
  output wire         pipe_tx2_compliance_o    ,
  output wire [ 1:0]  pipe_tx2_char_is_k_o     ,
  output wire [15:0]  pipe_tx2_data_o          ,
  output wire         pipe_tx2_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx2_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 3
  output  wire [ 1:0] pipe_rx3_char_is_k_o     ,
  output  wire [15:0] pipe_rx3_data_o         ,
  output  wire        pipe_rx3_valid_o         ,
  output  wire        pipe_rx3_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx3_status_o        ,
  output  wire        pipe_rx3_phy_status_o    ,
  output  wire        pipe_rx3_elec_idle_o     ,
  input   wire        pipe_rx3_polarity_i      ,
  input   wire        pipe_tx3_compliance_i    ,
  input   wire [ 1:0] pipe_tx3_char_is_k_i     ,
  input   wire [15:0] pipe_tx3_data_i          ,
  input   wire        pipe_tx3_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx3_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx3_char_is_k_i     ,
  input  wire [15:0]  pipe_rx3_data_i         ,
  input  wire         pipe_rx3_valid_i         ,
  input  wire         pipe_rx3_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx3_status_i        ,
  input  wire         pipe_rx3_phy_status_i    ,
  input  wire         pipe_rx3_elec_idle_i     ,
  output wire         pipe_rx3_polarity_o      ,
  output wire         pipe_tx3_compliance_o    ,
  output wire [ 1:0]  pipe_tx3_char_is_k_o     ,
  output wire [15:0]  pipe_tx3_data_o          ,
  output wire         pipe_tx3_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx3_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 4
  output  wire [ 1:0] pipe_rx4_char_is_k_o     ,
  output  wire [15:0] pipe_rx4_data_o         ,
  output  wire        pipe_rx4_valid_o         ,
  output  wire        pipe_rx4_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx4_status_o        ,
  output  wire        pipe_rx4_phy_status_o    ,
  output  wire        pipe_rx4_elec_idle_o     ,
  input   wire        pipe_rx4_polarity_i      ,
  input   wire        pipe_tx4_compliance_i    ,
  input   wire [ 1:0] pipe_tx4_char_is_k_i     ,
  input   wire [15:0] pipe_tx4_data_i          ,
  input   wire        pipe_tx4_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx4_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx4_char_is_k_i     ,
  input  wire [15:0]  pipe_rx4_data_i         ,
  input  wire         pipe_rx4_valid_i         ,
  input  wire         pipe_rx4_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx4_status_i        ,
  input  wire         pipe_rx4_phy_status_i    ,
  input  wire         pipe_rx4_elec_idle_i     ,
  output wire         pipe_rx4_polarity_o      ,
  output wire         pipe_tx4_compliance_o    ,
  output wire [ 1:0]  pipe_tx4_char_is_k_o     ,
  output wire [15:0]  pipe_tx4_data_o          ,
  output wire         pipe_tx4_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx4_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 5
  output  wire [ 1:0] pipe_rx5_char_is_k_o     ,
  output  wire [15:0] pipe_rx5_data_o         ,
  output  wire        pipe_rx5_valid_o         ,
  output  wire        pipe_rx5_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx5_status_o        ,
  output  wire        pipe_rx5_phy_status_o    ,
  output  wire        pipe_rx5_elec_idle_o     ,
  input   wire        pipe_rx5_polarity_i      ,
  input   wire        pipe_tx5_compliance_i    ,
  input   wire [ 1:0] pipe_tx5_char_is_k_i     ,
  input   wire [15:0] pipe_tx5_data_i          ,
  input   wire        pipe_tx5_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx5_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx5_char_is_k_i     ,
  input  wire [15:0]  pipe_rx5_data_i         ,
  input  wire         pipe_rx5_valid_i         ,
  input  wire         pipe_rx5_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx5_status_i        ,
  input  wire         pipe_rx5_phy_status_i    ,
  input  wire         pipe_rx5_elec_idle_i     ,
  output wire         pipe_rx5_polarity_o      ,
  output wire         pipe_tx5_compliance_o    ,
  output wire [ 1:0]  pipe_tx5_char_is_k_o     ,
  output wire [15:0]  pipe_tx5_data_o          ,
  output wire         pipe_tx5_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx5_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 6
  output  wire [ 1:0] pipe_rx6_char_is_k_o     ,
  output  wire [15:0] pipe_rx6_data_o         ,
  output  wire        pipe_rx6_valid_o         ,
  output  wire        pipe_rx6_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx6_status_o        ,
  output  wire        pipe_rx6_phy_status_o    ,
  output  wire        pipe_rx6_elec_idle_o     ,
  input   wire        pipe_rx6_polarity_i      ,
  input   wire        pipe_tx6_compliance_i    ,
  input   wire [ 1:0] pipe_tx6_char_is_k_i     ,
  input   wire [15:0] pipe_tx6_data_i          ,
  input   wire        pipe_tx6_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx6_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx6_char_is_k_i     ,
  input  wire [15:0]  pipe_rx6_data_i         ,
  input  wire         pipe_rx6_valid_i         ,
  input  wire         pipe_rx6_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx6_status_i        ,
  input  wire         pipe_rx6_phy_status_i    ,
  input  wire         pipe_rx6_elec_idle_i     ,
  output wire         pipe_rx6_polarity_o      ,
  output wire         pipe_tx6_compliance_o    ,
  output wire [ 1:0]  pipe_tx6_char_is_k_o     ,
  output wire [15:0]  pipe_tx6_data_o          ,
  output wire         pipe_tx6_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx6_powerdown_o     ,

  // Pipe Per-Lane Signals - Lane 7
  output  wire [ 1:0] pipe_rx7_char_is_k_o     ,
  output  wire [15:0] pipe_rx7_data_o         ,
  output  wire        pipe_rx7_valid_o         ,
  output  wire        pipe_rx7_chanisaligned_o ,
  output  wire [ 2:0] pipe_rx7_status_o        ,
  output  wire        pipe_rx7_phy_status_o    ,
  output  wire        pipe_rx7_elec_idle_o     ,
  input   wire        pipe_rx7_polarity_i      ,
  input   wire        pipe_tx7_compliance_i    ,
  input   wire [ 1:0] pipe_tx7_char_is_k_i     ,
  input   wire [15:0] pipe_tx7_data_i          ,
  input   wire        pipe_tx7_elec_idle_i     ,
  input   wire [ 1:0] pipe_tx7_powerdown_i     ,

  input  wire [ 1:0]  pipe_rx7_char_is_k_i     ,
  input  wire [15:0]  pipe_rx7_data_i         ,
  input  wire         pipe_rx7_valid_i         ,
  input  wire         pipe_rx7_chanisaligned_i ,
  input  wire [ 2:0]  pipe_rx7_status_i        ,
  input  wire         pipe_rx7_phy_status_i    ,
  input  wire         pipe_rx7_elec_idle_i     ,
  output wire         pipe_rx7_polarity_o      ,
  output wire         pipe_tx7_compliance_o    ,
  output wire [ 1:0]  pipe_tx7_char_is_k_o     ,
  output wire [15:0]  pipe_tx7_data_o          ,
  output wire         pipe_tx7_elec_idle_o     ,
  output wire [ 1:0]  pipe_tx7_powerdown_o     ,

  // Non PIPE signals
  input   wire        pipe_clk               ,
  input   wire        rst_n
);

  //******************************************************************//
  // Reality check.                                                   //
  //******************************************************************//
  
  //synthesis translate_off
  //   initial begin
  //      $display("[%t] %m LINK_CAP_MAX_LINK_WIDTH %0d  PIPE_PIPELINE_STAGES %0d", 
  //                 $time, LINK_CAP_MAX_LINK_WIDTH, PIPE_PIPELINE_STAGES);
  //   end
  //synthesis translate_on

  generate

model_ap2_tst_pcie_pipe_misc # (

      .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

    )
    model_ap2_tst_pipe_misc_i (

      .pipe_tx_rcvr_det_i(pipe_tx_rcvr_det_i),
      .pipe_tx_reset_i(pipe_tx_reset_i),
      .pipe_tx_rate_i(pipe_tx_rate_i),
      .pipe_tx_deemph_i(pipe_tx_deemph_i),
      .pipe_tx_margin_i(pipe_tx_margin_i),
      .pipe_tx_swing_i(pipe_tx_swing_i),

      .pipe_tx_rcvr_det_o(pipe_tx_rcvr_det_o),
      .pipe_tx_reset_o(pipe_tx_reset_o),
      .pipe_tx_rate_o(pipe_tx_rate_o),
      .pipe_tx_deemph_o(pipe_tx_deemph_o),
      .pipe_tx_margin_o(pipe_tx_margin_o),
      .pipe_tx_swing_o(pipe_tx_swing_o)          ,

      .pipe_clk(pipe_clk),
      .rst_n(rst_n)
  );


model_ap2_tst_pcie_pipe_lane # (

      .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

    )
    model_ap2_tst_pipe_lane_0_i (

      .pipe_rx_char_is_k_o(pipe_rx0_char_is_k_o),
      .pipe_rx_data_o(pipe_rx0_data_o),
      .pipe_rx_valid_o(pipe_rx0_valid_o),
      .pipe_rx_chanisaligned_o(pipe_rx0_chanisaligned_o),
      .pipe_rx_status_o(pipe_rx0_status_o),
      .pipe_rx_phy_status_o(pipe_rx0_phy_status_o),
      .pipe_rx_elec_idle_o(pipe_rx0_elec_idle_o),
      .pipe_rx_polarity_i(pipe_rx0_polarity_i),
      .pipe_tx_compliance_i(pipe_tx0_compliance_i),
      .pipe_tx_char_is_k_i(pipe_tx0_char_is_k_i),
      .pipe_tx_data_i(pipe_tx0_data_i),
      .pipe_tx_elec_idle_i(pipe_tx0_elec_idle_i),
      .pipe_tx_powerdown_i(pipe_tx0_powerdown_i),

      .pipe_rx_char_is_k_i(pipe_rx0_char_is_k_i),
      .pipe_rx_data_i(pipe_rx0_data_i),
      .pipe_rx_valid_i(pipe_rx0_valid_i),
      .pipe_rx_chanisaligned_i(pipe_rx0_chanisaligned_i),
      .pipe_rx_status_i(pipe_rx0_status_i),
      .pipe_rx_phy_status_i(pipe_rx0_phy_status_i),
      .pipe_rx_elec_idle_i(pipe_rx0_elec_idle_i),
      .pipe_rx_polarity_o(pipe_rx0_polarity_o),
      .pipe_tx_compliance_o(pipe_tx0_compliance_o),
      .pipe_tx_char_is_k_o(pipe_tx0_char_is_k_o),
      .pipe_tx_data_o(pipe_tx0_data_o),
      .pipe_tx_elec_idle_o(pipe_tx0_elec_idle_o),
      .pipe_tx_powerdown_o(pipe_tx0_powerdown_o),

      .pipe_clk(pipe_clk),
      .rst_n(rst_n)

    );

    if (LINK_CAP_MAX_LINK_WIDTH >= 2) begin : pipe_2_lane

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_1_i (

        .pipe_rx_char_is_k_o(pipe_rx1_char_is_k_o),
        .pipe_rx_data_o(pipe_rx1_data_o),
        .pipe_rx_valid_o(pipe_rx1_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx1_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx1_status_o),
        .pipe_rx_phy_status_o(pipe_rx1_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx1_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx1_polarity_i),
        .pipe_tx_compliance_i(pipe_tx1_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx1_char_is_k_i),
        .pipe_tx_data_i(pipe_tx1_data_i),
        .pipe_tx_elec_idle_i(pipe_tx1_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx1_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx1_char_is_k_i),
        .pipe_rx_data_i(pipe_rx1_data_i),
        .pipe_rx_valid_i(pipe_rx1_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx1_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx1_status_i),
        .pipe_rx_phy_status_i(pipe_rx1_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx1_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx1_polarity_o),
        .pipe_tx_compliance_o(pipe_tx1_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx1_char_is_k_o),
        .pipe_tx_data_o(pipe_tx1_data_o),
        .pipe_tx_elec_idle_o(pipe_tx1_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx1_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

    end // if (LINK_CAP_MAX_LINK_WIDTH >= 2)
    else
    begin
      assign pipe_rx1_char_is_k_o = 2'b00;
      assign pipe_rx1_data_o = 16'h0000;
      assign pipe_rx1_valid_o = 1'b0;
      assign pipe_rx1_chanisaligned_o = 1'b0;
      assign pipe_rx1_status_o = 3'b000;
      assign pipe_rx1_phy_status_o = 1'b0;
      assign pipe_rx1_elec_idle_o = 1'b1;
      assign pipe_rx1_polarity_o = 1'b0;
      assign pipe_tx1_compliance_o = 1'b0;
      assign pipe_tx1_char_is_k_o = 2'b00;
      assign pipe_tx1_data_o = 16'h0000;
      assign pipe_tx1_elec_idle_o = 1'b1;
      assign pipe_tx1_powerdown_o = 2'b00;
    end // if !(LINK_CAP_MAX_LINK_WIDTH >= 2)

    if (LINK_CAP_MAX_LINK_WIDTH >= 4) begin : pipe_4_lane

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)
      )
      model_ap2_tst_pipe_lane_2_i (

        .pipe_rx_char_is_k_o(pipe_rx2_char_is_k_o),
        .pipe_rx_data_o(pipe_rx2_data_o),
        .pipe_rx_valid_o(pipe_rx2_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx2_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx2_status_o),
        .pipe_rx_phy_status_o(pipe_rx2_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx2_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx2_polarity_i),
        .pipe_tx_compliance_i(pipe_tx2_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx2_char_is_k_i),
        .pipe_tx_data_i(pipe_tx2_data_i),
        .pipe_tx_elec_idle_i(pipe_tx2_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx2_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx2_char_is_k_i),
        .pipe_rx_data_i(pipe_rx2_data_i),
        .pipe_rx_valid_i(pipe_rx2_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx2_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx2_status_i),
        .pipe_rx_phy_status_i(pipe_rx2_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx2_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx2_polarity_o),
        .pipe_tx_compliance_o(pipe_tx2_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx2_char_is_k_o),
        .pipe_tx_data_o(pipe_tx2_data_o),
        .pipe_tx_elec_idle_o(pipe_tx2_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx2_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_3_i (

        .pipe_rx_char_is_k_o(pipe_rx3_char_is_k_o),
        .pipe_rx_data_o(pipe_rx3_data_o),
        .pipe_rx_valid_o(pipe_rx3_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx3_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx3_status_o),
        .pipe_rx_phy_status_o(pipe_rx3_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx3_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx3_polarity_i),
        .pipe_tx_compliance_i(pipe_tx3_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx3_char_is_k_i),
        .pipe_tx_data_i(pipe_tx3_data_i),
        .pipe_tx_elec_idle_i(pipe_tx3_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx3_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx3_char_is_k_i),
        .pipe_rx_data_i(pipe_rx3_data_i),
        .pipe_rx_valid_i(pipe_rx3_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx3_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx3_status_i),
        .pipe_rx_phy_status_i(pipe_rx3_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx3_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx3_polarity_o),
        .pipe_tx_compliance_o(pipe_tx3_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx3_char_is_k_o),
        .pipe_tx_data_o(pipe_tx3_data_o),
        .pipe_tx_elec_idle_o(pipe_tx3_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx3_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

    end // if (LINK_CAP_MAX_LINK_WIDTH >= 4)
    else
    begin
      assign pipe_rx2_char_is_k_o = 2'b00;
      assign pipe_rx2_data_o = 16'h0000;
      assign pipe_rx2_valid_o = 1'b0;
      assign pipe_rx2_chanisaligned_o = 1'b0;
      assign pipe_rx2_status_o = 3'b000;
      assign pipe_rx2_phy_status_o = 1'b0;
      assign pipe_rx2_elec_idle_o = 1'b1;
      assign pipe_rx2_polarity_o = 1'b0;
      assign pipe_tx2_compliance_o = 1'b0;
      assign pipe_tx2_char_is_k_o = 2'b00;
      assign pipe_tx2_data_o = 16'h0000;
      assign pipe_tx2_elec_idle_o = 1'b1;
      assign pipe_tx2_powerdown_o = 2'b00;

      assign pipe_rx3_char_is_k_o = 2'b00;
      assign pipe_rx3_data_o = 16'h0000;
      assign pipe_rx3_valid_o = 1'b0;
      assign pipe_rx3_chanisaligned_o = 1'b0;
      assign pipe_rx3_status_o = 3'b000;
      assign pipe_rx3_phy_status_o = 1'b0;
      assign pipe_rx3_elec_idle_o = 1'b1;
      assign pipe_rx3_polarity_o = 1'b0;
      assign pipe_tx3_compliance_o = 1'b0;
      assign pipe_tx3_char_is_k_o = 2'b00;
      assign pipe_tx3_data_o = 16'h0000;
      assign pipe_tx3_elec_idle_o = 1'b1;
      assign pipe_tx3_powerdown_o = 2'b00;
    end // if !(LINK_CAP_MAX_LINK_WIDTH >= 4)

    if (LINK_CAP_MAX_LINK_WIDTH >= 8) begin : pipe_8_lane

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_4_i (

        .pipe_rx_char_is_k_o(pipe_rx4_char_is_k_o),
        .pipe_rx_data_o(pipe_rx4_data_o),
        .pipe_rx_valid_o(pipe_rx4_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx4_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx4_status_o),
        .pipe_rx_phy_status_o(pipe_rx4_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx4_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx4_polarity_i),
        .pipe_tx_compliance_i(pipe_tx4_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx4_char_is_k_i),
        .pipe_tx_data_i(pipe_tx4_data_i),
        .pipe_tx_elec_idle_i(pipe_tx4_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx4_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx4_char_is_k_i),
        .pipe_rx_data_i(pipe_rx4_data_i),
        .pipe_rx_valid_i(pipe_rx4_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx4_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx4_status_i),
        .pipe_rx_phy_status_i(pipe_rx4_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx4_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx4_polarity_o),
        .pipe_tx_compliance_o(pipe_tx4_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx4_char_is_k_o),
        .pipe_tx_data_o(pipe_tx4_data_o),
        .pipe_tx_elec_idle_o(pipe_tx4_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx4_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_5_i (

        .pipe_rx_char_is_k_o(pipe_rx5_char_is_k_o),
        .pipe_rx_data_o(pipe_rx5_data_o),
        .pipe_rx_valid_o(pipe_rx5_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx5_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx5_status_o),
        .pipe_rx_phy_status_o(pipe_rx5_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx5_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx5_polarity_i),
        .pipe_tx_compliance_i(pipe_tx5_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx5_char_is_k_i),
        .pipe_tx_data_i(pipe_tx5_data_i),
        .pipe_tx_elec_idle_i(pipe_tx5_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx5_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx5_char_is_k_i),
        .pipe_rx_data_i(pipe_rx5_data_i),
        .pipe_rx_valid_i(pipe_rx5_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx5_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx5_status_i),
        .pipe_rx_phy_status_i(pipe_rx5_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx5_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx5_polarity_o),
        .pipe_tx_compliance_o(pipe_tx5_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx5_char_is_k_o),
        .pipe_tx_data_o(pipe_tx5_data_o),
        .pipe_tx_elec_idle_o(pipe_tx5_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx5_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_6_i (

        .pipe_rx_char_is_k_o(pipe_rx6_char_is_k_o),
        .pipe_rx_data_o(pipe_rx6_data_o),
        .pipe_rx_valid_o(pipe_rx6_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx6_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx6_status_o),
        .pipe_rx_phy_status_o(pipe_rx6_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx6_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx6_polarity_i),
        .pipe_tx_compliance_i(pipe_tx6_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx6_char_is_k_i),
        .pipe_tx_data_i(pipe_tx6_data_i),
        .pipe_tx_elec_idle_i(pipe_tx6_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx6_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx6_char_is_k_i),
        .pipe_rx_data_i(pipe_rx6_data_i),
        .pipe_rx_valid_i(pipe_rx6_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx6_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx6_status_i),
        .pipe_rx_phy_status_i(pipe_rx6_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx6_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx6_polarity_o),
        .pipe_tx_compliance_o(pipe_tx6_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx6_char_is_k_o),
        .pipe_tx_data_o(pipe_tx6_data_o),
        .pipe_tx_elec_idle_o(pipe_tx6_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx6_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

model_ap2_tst_pcie_pipe_lane # (

        .PIPE_PIPELINE_STAGES(PIPE_PIPELINE_STAGES)

      )
      model_ap2_tst_pipe_lane_7_i (

        .pipe_rx_char_is_k_o(pipe_rx7_char_is_k_o),
        .pipe_rx_data_o(pipe_rx7_data_o),
        .pipe_rx_valid_o(pipe_rx7_valid_o),
        .pipe_rx_chanisaligned_o(pipe_rx7_chanisaligned_o),
        .pipe_rx_status_o(pipe_rx7_status_o),
        .pipe_rx_phy_status_o(pipe_rx7_phy_status_o),
        .pipe_rx_elec_idle_o(pipe_rx7_elec_idle_o),
        .pipe_rx_polarity_i(pipe_rx7_polarity_i),
        .pipe_tx_compliance_i(pipe_tx7_compliance_i),
        .pipe_tx_char_is_k_i(pipe_tx7_char_is_k_i),
        .pipe_tx_data_i(pipe_tx7_data_i),
        .pipe_tx_elec_idle_i(pipe_tx7_elec_idle_i),
        .pipe_tx_powerdown_i(pipe_tx7_powerdown_i),

        .pipe_rx_char_is_k_i(pipe_rx7_char_is_k_i),
        .pipe_rx_data_i(pipe_rx7_data_i),
        .pipe_rx_valid_i(pipe_rx7_valid_i),
        .pipe_rx_chanisaligned_i(pipe_rx7_chanisaligned_i),
        .pipe_rx_status_i(pipe_rx7_status_i),
        .pipe_rx_phy_status_i(pipe_rx7_phy_status_i),
        .pipe_rx_elec_idle_i(pipe_rx7_elec_idle_i),
        .pipe_rx_polarity_o(pipe_rx7_polarity_o),
        .pipe_tx_compliance_o(pipe_tx7_compliance_o),
        .pipe_tx_char_is_k_o(pipe_tx7_char_is_k_o),
        .pipe_tx_data_o(pipe_tx7_data_o),
        .pipe_tx_elec_idle_o(pipe_tx7_elec_idle_o),
        .pipe_tx_powerdown_o(pipe_tx7_powerdown_o),

        .pipe_clk(pipe_clk),
        .rst_n(rst_n)

      );

    end // if (LINK_CAP_MAX_LINK_WIDTH >= 8)
    else
    begin
      assign pipe_rx4_char_is_k_o = 2'b00;
      assign pipe_rx4_data_o = 16'h0000;
      assign pipe_rx4_valid_o = 1'b0;
      assign pipe_rx4_chanisaligned_o = 1'b0;
      assign pipe_rx4_status_o = 3'b000;
      assign pipe_rx4_phy_status_o = 1'b0;
      assign pipe_rx4_elec_idle_o = 1'b1;
      assign pipe_rx4_polarity_o = 1'b0;
      assign pipe_tx4_compliance_o = 1'b0;
      assign pipe_tx4_char_is_k_o = 2'b00;
      assign pipe_tx4_data_o = 16'h0000;
      assign pipe_tx4_elec_idle_o = 1'b1;
      assign pipe_tx4_powerdown_o = 2'b00;

      assign pipe_rx5_char_is_k_o = 2'b00;
      assign pipe_rx5_data_o = 16'h0000;
      assign pipe_rx5_valid_o = 1'b0;
      assign pipe_rx5_chanisaligned_o = 1'b0;
      assign pipe_rx5_status_o = 3'b000;
      assign pipe_rx5_phy_status_o = 1'b0;
      assign pipe_rx5_elec_idle_o = 1'b1;
      assign pipe_rx5_polarity_o = 1'b0;
      assign pipe_tx5_compliance_o = 1'b0;
      assign pipe_tx5_char_is_k_o = 2'b00;
      assign pipe_tx5_data_o = 16'h0000;
      assign pipe_tx5_elec_idle_o = 1'b1;
      assign pipe_tx5_powerdown_o = 2'b00;

      assign pipe_rx6_char_is_k_o = 2'b00;
      assign pipe_rx6_data_o = 16'h0000;
      assign pipe_rx6_valid_o = 1'b0;
      assign pipe_rx6_chanisaligned_o = 1'b0;
      assign pipe_rx6_status_o = 3'b000;
      assign pipe_rx6_phy_status_o = 1'b0;
      assign pipe_rx6_elec_idle_o = 1'b1;
      assign pipe_rx6_polarity_o = 1'b0;
      assign pipe_tx6_compliance_o = 1'b0;
      assign pipe_tx6_char_is_k_o = 2'b00;
      assign pipe_tx6_data_o = 16'h0000;
      assign pipe_tx6_elec_idle_o = 1'b1;
      assign pipe_tx6_powerdown_o = 2'b00;

      assign pipe_rx7_char_is_k_o = 2'b00;
      assign pipe_rx7_data_o = 16'h0000;
      assign pipe_rx7_valid_o = 1'b0;
      assign pipe_rx7_chanisaligned_o = 1'b0;
      assign pipe_rx7_status_o = 3'b000;
      assign pipe_rx7_phy_status_o = 1'b0;
      assign pipe_rx7_elec_idle_o = 1'b1;
      assign pipe_rx7_polarity_o = 1'b0;
      assign pipe_tx7_compliance_o = 1'b0;
      assign pipe_tx7_char_is_k_o = 2'b00;
      assign pipe_tx7_data_o = 16'h0000;
      assign pipe_tx7_elec_idle_o = 1'b1;
      assign pipe_tx7_powerdown_o = 2'b00;
    end // if !(LINK_CAP_MAX_LINK_WIDTH >= 8)

  endgenerate

endmodule



`timescale 1ns/1ps
module model_ap2_tst_pcie_pipe_misc #
(
    parameter        PIPE_PIPELINE_STAGES = 0,    // 0 - 0 stages, 1 - 1 stage, 2 - 2 stages
    parameter TCQ  = 1 // synthesis warning solved: parameter declaration becomes local
)
(

    input   wire        pipe_tx_rcvr_det_i       ,     // PIPE Tx Receiver Detect
    input   wire        pipe_tx_reset_i          ,     // PIPE Tx Reset
    input   wire        pipe_tx_rate_i           ,     // PIPE Tx Rate
    input   wire        pipe_tx_deemph_i         ,     // PIPE Tx Deemphasis
    input   wire [2:0]  pipe_tx_margin_i         ,     // PIPE Tx Margin
    input   wire        pipe_tx_swing_i          ,     // PIPE Tx Swing

    output  wire        pipe_tx_rcvr_det_o       ,     // Pipelined PIPE Tx Receiver Detect
    output  wire        pipe_tx_reset_o          ,     // Pipelined PIPE Tx Reset
    output  wire        pipe_tx_rate_o           ,     // Pipelined PIPE Tx Rate
    output  wire        pipe_tx_deemph_o         ,     // Pipelined PIPE Tx Deemphasis
    output  wire [2:0]  pipe_tx_margin_o         ,     // Pipelined PIPE Tx Margin
    output  wire        pipe_tx_swing_o          ,     // Pipelined PIPE Tx Swing

    input   wire        pipe_clk                ,      // PIPE Clock
    input   wire        rst_n                          // Reset
);

//******************************************************************//
// Reality check.                                                   //
//******************************************************************//

//    parameter TCQ  = 1;      // clock to out delay model

    generate

    if (PIPE_PIPELINE_STAGES == 0) begin : pipe_stages_0

        assign pipe_tx_rcvr_det_o = pipe_tx_rcvr_det_i;
        assign pipe_tx_reset_o  = pipe_tx_reset_i;
        assign pipe_tx_rate_o = pipe_tx_rate_i;
        assign pipe_tx_deemph_o = pipe_tx_deemph_i;
        assign pipe_tx_margin_o = pipe_tx_margin_i;
        assign pipe_tx_swing_o = pipe_tx_swing_i;

    end // if (PIPE_PIPELINE_STAGES == 0)
    else if (PIPE_PIPELINE_STAGES == 1) begin : pipe_stages_1

    reg                pipe_tx_rcvr_det_q       ;
    reg                pipe_tx_reset_q          ;
    reg                pipe_tx_rate_q           ;
    reg                pipe_tx_deemph_q         ;
    reg [2:0]          pipe_tx_margin_q         ;
    reg                pipe_tx_swing_q          ;

        always @(posedge pipe_clk) begin

        if (rst_n)
        begin

            pipe_tx_rcvr_det_q <= #TCQ 0;
            pipe_tx_reset_q  <= #TCQ 1'b1;
            pipe_tx_rate_q <= #TCQ 0;
            pipe_tx_deemph_q <= #TCQ 1'b1;
            pipe_tx_margin_q <= #TCQ 0;
            pipe_tx_swing_q <= #TCQ 0;

        end
        else
        begin

            pipe_tx_rcvr_det_q <= #TCQ pipe_tx_rcvr_det_i;
            pipe_tx_reset_q  <= #TCQ pipe_tx_reset_i;
            pipe_tx_rate_q <= #TCQ pipe_tx_rate_i;
            pipe_tx_deemph_q <= #TCQ pipe_tx_deemph_i;
            pipe_tx_margin_q <= #TCQ pipe_tx_margin_i;
            pipe_tx_swing_q <= #TCQ pipe_tx_swing_i;

          end

        end

        assign pipe_tx_rcvr_det_o = pipe_tx_rcvr_det_q;
        assign pipe_tx_reset_o  = pipe_tx_reset_q;
        assign pipe_tx_rate_o = pipe_tx_rate_q;
        assign pipe_tx_deemph_o = pipe_tx_deemph_q;
        assign pipe_tx_margin_o = pipe_tx_margin_q;
        assign pipe_tx_swing_o = pipe_tx_swing_q;

    end // if (PIPE_PIPELINE_STAGES == 1)
    else if (PIPE_PIPELINE_STAGES == 2) begin : pipe_stages_2

    reg                pipe_tx_rcvr_det_q       ;
    reg                pipe_tx_reset_q          ;
    reg                pipe_tx_rate_q           ;
    reg                pipe_tx_deemph_q         ;
    reg [2:0]          pipe_tx_margin_q         ;
    reg                pipe_tx_swing_q          ;

    reg                pipe_tx_rcvr_det_qq      ;
    reg                pipe_tx_reset_qq         ;
    reg                pipe_tx_rate_qq          ;
    reg                pipe_tx_deemph_qq        ;
    reg [2:0]          pipe_tx_margin_qq        ;
    reg                pipe_tx_swing_qq         ;

        always @(posedge pipe_clk) begin

        if (rst_n)
        begin

            pipe_tx_rcvr_det_q <= #TCQ 0;
            pipe_tx_reset_q  <= #TCQ 1'b1;
            pipe_tx_rate_q <= #TCQ 0;
            pipe_tx_deemph_q <= #TCQ 1'b1;
            pipe_tx_margin_q <= #TCQ 0;
            pipe_tx_swing_q <= #TCQ 0;

            pipe_tx_rcvr_det_qq <= #TCQ 0;
            pipe_tx_reset_qq  <= #TCQ 1'b1;
            pipe_tx_rate_qq <= #TCQ 0;
            pipe_tx_deemph_qq <= #TCQ 1'b1;
            pipe_tx_margin_qq <= #TCQ 0;
            pipe_tx_swing_qq <= #TCQ 0;

        end
        else
        begin

            pipe_tx_rcvr_det_q <= #TCQ pipe_tx_rcvr_det_i;
            pipe_tx_reset_q  <= #TCQ pipe_tx_reset_i;
            pipe_tx_rate_q <= #TCQ pipe_tx_rate_i;
            pipe_tx_deemph_q <= #TCQ pipe_tx_deemph_i;
            pipe_tx_margin_q <= #TCQ pipe_tx_margin_i;
            pipe_tx_swing_q <= #TCQ pipe_tx_swing_i;

            pipe_tx_rcvr_det_qq <= #TCQ pipe_tx_rcvr_det_q;
            pipe_tx_reset_qq  <= #TCQ pipe_tx_reset_q;
            pipe_tx_rate_qq <= #TCQ pipe_tx_rate_q;
            pipe_tx_deemph_qq <= #TCQ pipe_tx_deemph_q;
            pipe_tx_margin_qq <= #TCQ pipe_tx_margin_q;
            pipe_tx_swing_qq <= #TCQ pipe_tx_swing_q;

          end

        end

        assign pipe_tx_rcvr_det_o = pipe_tx_rcvr_det_qq;
        assign pipe_tx_reset_o  = pipe_tx_reset_qq;
        assign pipe_tx_rate_o = pipe_tx_rate_qq;
        assign pipe_tx_deemph_o = pipe_tx_deemph_qq;
        assign pipe_tx_margin_o = pipe_tx_margin_qq;
        assign pipe_tx_swing_o = pipe_tx_swing_qq;

    end // if (PIPE_PIPELINE_STAGES == 2)

    endgenerate

endmodule



`timescale 1ns/1ps
module model_ap2_tst_pcie_pipe_lane #
(
    parameter        PIPE_PIPELINE_STAGES = 0,    // 0 - 0 stages, 1 - 1 stage, 2 - 2 stages
    parameter TCQ  = 1 // synthesis warning solved : parameter declaration becomes local
)
(
    output  wire [ 1:0] pipe_rx_char_is_k_o     ,    // Pipelined PIPE Rx Char Is K
    output  wire [15:0] pipe_rx_data_o          ,    // Pipelined PIPE Rx Data
    output  wire        pipe_rx_valid_o         ,    // Pipelined PIPE Rx Data Valid
    output  wire        pipe_rx_chanisaligned_o ,    // Pipelined PIPE Rx Chan Is Aligned
    output  wire [ 2:0] pipe_rx_status_o        ,    // Pipelined PIPE Rx Status
    output  wire        pipe_rx_phy_status_o    ,    // Pipelined PIPE Rx Phy Status
    output  wire        pipe_rx_elec_idle_o     ,    // Pipelined PIPE Rx Electrical Idle
    input   wire        pipe_rx_polarity_i      ,    // PIPE Rx Polarity
    input   wire        pipe_tx_compliance_i    ,    // PIPE Tx Compliance
    input   wire [ 1:0] pipe_tx_char_is_k_i     ,    // PIPE Tx Char Is K
    input   wire [15:0] pipe_tx_data_i          ,    // PIPE Tx Data
    input   wire        pipe_tx_elec_idle_i     ,    // PIPE Tx Electrical Idle
    input   wire [ 1:0] pipe_tx_powerdown_i     ,    // PIPE Tx Powerdown

    input  wire [ 1:0]  pipe_rx_char_is_k_i     ,    // PIPE Rx Char Is K
    input  wire [15:0]  pipe_rx_data_i          ,    // PIPE Rx Data
    input  wire         pipe_rx_valid_i         ,    // PIPE Rx Data Valid
    input  wire         pipe_rx_chanisaligned_i ,    // PIPE Rx Chan Is Aligned
    input  wire [ 2:0]  pipe_rx_status_i        ,    // PIPE Rx Status
    input  wire         pipe_rx_phy_status_i    ,    // PIPE Rx Phy Status
    input  wire         pipe_rx_elec_idle_i     ,    // PIPE Rx Electrical Idle
    output wire         pipe_rx_polarity_o      ,    // Pipelined PIPE Rx Polarity
    output wire         pipe_tx_compliance_o    ,    // Pipelined PIPE Tx Compliance
    output wire [ 1:0]  pipe_tx_char_is_k_o     ,    // Pipelined PIPE Tx Char Is K
    output wire [15:0]  pipe_tx_data_o          ,    // Pipelined PIPE Tx Data
    output wire         pipe_tx_elec_idle_o     ,    // Pipelined PIPE Tx Electrical Idle
    output wire [ 1:0]  pipe_tx_powerdown_o     ,    // Pipelined PIPE Tx Powerdown

    input   wire        pipe_clk                ,    // PIPE Clock
    input   wire        rst_n                        // Reset
);

  //******************************************************************//
  // Reality check.                                                   //
  //******************************************************************//

//    parameter TCQ  = 1;      // clock to out delay model

    generate

    if (PIPE_PIPELINE_STAGES == 0) begin : pipe_stages_0

        assign pipe_rx_char_is_k_o = pipe_rx_char_is_k_i;
        assign pipe_rx_data_o = pipe_rx_data_i;
        assign pipe_rx_valid_o = pipe_rx_valid_i;
        assign pipe_rx_chanisaligned_o = pipe_rx_chanisaligned_i;
        assign pipe_rx_status_o = pipe_rx_status_i;
        assign pipe_rx_phy_status_o = pipe_rx_phy_status_i;
        assign pipe_rx_elec_idle_o = pipe_rx_elec_idle_i;

        assign pipe_rx_polarity_o = pipe_rx_polarity_i;
        assign pipe_tx_compliance_o = pipe_tx_compliance_i;
        assign pipe_tx_char_is_k_o = pipe_tx_char_is_k_i;
        assign pipe_tx_data_o = pipe_tx_data_i;
        assign pipe_tx_elec_idle_o = pipe_tx_elec_idle_i;
        assign pipe_tx_powerdown_o = pipe_tx_powerdown_i;

    end // if (PIPE_PIPELINE_STAGES == 0)
    else if (PIPE_PIPELINE_STAGES == 1) begin : pipe_stages_1

    reg [ 1:0]          pipe_rx_char_is_k_q     ;
    reg [15:0]          pipe_rx_data_q          ;
    reg                 pipe_rx_valid_q         ;
    reg                 pipe_rx_chanisaligned_q ;
    reg [ 2:0]          pipe_rx_status_q        ;
    reg                 pipe_rx_phy_status_q    ;
    reg                 pipe_rx_elec_idle_q     ;

    reg                 pipe_rx_polarity_q      ;
    reg                 pipe_tx_compliance_q    ;
    reg [ 1:0]          pipe_tx_char_is_k_q     ;
    reg [15:0]          pipe_tx_data_q          ;
    reg                 pipe_tx_elec_idle_q     ;
    reg [ 1:0]          pipe_tx_powerdown_q     ;

        always @(posedge pipe_clk) begin

        if (rst_n) 
        begin

            pipe_rx_char_is_k_q <= #TCQ 0;
            pipe_rx_data_q <= #TCQ 0;
            pipe_rx_valid_q <= #TCQ 0;
            pipe_rx_chanisaligned_q <= #TCQ 0;
            pipe_rx_status_q <= #TCQ 0;
            pipe_rx_phy_status_q <= #TCQ 0;
            pipe_rx_elec_idle_q <= #TCQ 0;

            pipe_rx_polarity_q <= #TCQ 0;
            pipe_tx_compliance_q <= #TCQ 0;
            pipe_tx_char_is_k_q <= #TCQ 0;
            pipe_tx_data_q <= #TCQ 0;
            pipe_tx_elec_idle_q <= #TCQ 1'b1;
            pipe_tx_powerdown_q <= #TCQ 2'b10;

        end
        else 
        begin

            pipe_rx_char_is_k_q <= #TCQ pipe_rx_char_is_k_i;
            pipe_rx_data_q <= #TCQ pipe_rx_data_i;
            pipe_rx_valid_q <= #TCQ pipe_rx_valid_i;
            pipe_rx_chanisaligned_q <= #TCQ pipe_rx_chanisaligned_i;
            pipe_rx_status_q <= #TCQ pipe_rx_status_i;
            pipe_rx_phy_status_q <= #TCQ pipe_rx_phy_status_i;
            pipe_rx_elec_idle_q <= #TCQ pipe_rx_elec_idle_i;

            pipe_rx_polarity_q <= #TCQ pipe_rx_polarity_i;
            pipe_tx_compliance_q <= #TCQ pipe_tx_compliance_i;
            pipe_tx_char_is_k_q <= #TCQ pipe_tx_char_is_k_i;
            pipe_tx_data_q <= #TCQ pipe_tx_data_i;
            pipe_tx_elec_idle_q <= #TCQ pipe_tx_elec_idle_i;
            pipe_tx_powerdown_q <= #TCQ pipe_tx_powerdown_i;

          end

        end

        assign pipe_rx_char_is_k_o = pipe_rx_char_is_k_q;
        assign pipe_rx_data_o = pipe_rx_data_q;
        assign pipe_rx_valid_o = pipe_rx_valid_q;
        assign pipe_rx_chanisaligned_o = pipe_rx_chanisaligned_q;
        assign pipe_rx_status_o = pipe_rx_status_q;
        assign pipe_rx_phy_status_o = pipe_rx_phy_status_q;
        assign pipe_rx_elec_idle_o = pipe_rx_elec_idle_q;

        assign pipe_rx_polarity_o = pipe_rx_polarity_q;
        assign pipe_tx_compliance_o = pipe_tx_compliance_q;
        assign pipe_tx_char_is_k_o = pipe_tx_char_is_k_q;
        assign pipe_tx_data_o = pipe_tx_data_q;
        assign pipe_tx_elec_idle_o = pipe_tx_elec_idle_q;
        assign pipe_tx_powerdown_o = pipe_tx_powerdown_q;

    end // if (PIPE_PIPELINE_STAGES == 1)
    else if (PIPE_PIPELINE_STAGES == 2) begin : pipe_stages_2

    reg [ 1:0]          pipe_rx_char_is_k_q     ;
    reg [15:0]          pipe_rx_data_q          ;
    reg                 pipe_rx_valid_q         ;
    reg                 pipe_rx_chanisaligned_q ;
    reg [ 2:0]          pipe_rx_status_q        ;
    reg                 pipe_rx_phy_status_q    ;
    reg                 pipe_rx_elec_idle_q     ;

    reg                 pipe_rx_polarity_q      ;
    reg                 pipe_tx_compliance_q    ;
    reg [ 1:0]          pipe_tx_char_is_k_q     ;
    reg [15:0]          pipe_tx_data_q          ;
    reg                 pipe_tx_elec_idle_q     ;
    reg [ 1:0]          pipe_tx_powerdown_q     ;

    reg [ 1:0]          pipe_rx_char_is_k_qq    ;
    reg [15:0]          pipe_rx_data_qq         ;
    reg                 pipe_rx_valid_qq        ;
    reg                 pipe_rx_chanisaligned_qq;
    reg [ 2:0]          pipe_rx_status_qq       ;
    reg                 pipe_rx_phy_status_qq   ;
    reg                 pipe_rx_elec_idle_qq    ;

    reg                 pipe_rx_polarity_qq     ;
    reg                 pipe_tx_compliance_qq   ;
    reg [ 1:0]          pipe_tx_char_is_k_qq    ;
    reg [15:0]          pipe_tx_data_qq         ;
    reg                 pipe_tx_elec_idle_qq    ;
    reg [ 1:0]          pipe_tx_powerdown_qq    ;

        always @(posedge pipe_clk) begin

        if (rst_n) 
        begin

            pipe_rx_char_is_k_q <= #TCQ 0;
            pipe_rx_data_q <= #TCQ 0;
            pipe_rx_valid_q <= #TCQ 0;
            pipe_rx_chanisaligned_q <= #TCQ 0;
            pipe_rx_status_q <= #TCQ 0;
            pipe_rx_phy_status_q <= #TCQ 0;
            pipe_rx_elec_idle_q <= #TCQ 0;

            pipe_rx_polarity_q <= #TCQ 0;
            pipe_tx_compliance_q <= #TCQ 0;
            pipe_tx_char_is_k_q <= #TCQ 0;
            pipe_tx_data_q <= #TCQ 0;
            pipe_tx_elec_idle_q <= #TCQ 1'b1;
            pipe_tx_powerdown_q <= #TCQ 2'b10;

            pipe_rx_char_is_k_qq <= #TCQ 0;
            pipe_rx_data_qq <= #TCQ 0;
            pipe_rx_valid_qq <= #TCQ 0;
            pipe_rx_chanisaligned_qq <= #TCQ 0;
            pipe_rx_status_qq <= #TCQ 0;
            pipe_rx_phy_status_qq <= #TCQ 0;
            pipe_rx_elec_idle_qq <= #TCQ 0;

            pipe_rx_polarity_qq <= #TCQ 0;
            pipe_tx_compliance_qq <= #TCQ 0;
            pipe_tx_char_is_k_qq <= #TCQ 0;
            pipe_tx_data_qq <= #TCQ 0;
            pipe_tx_elec_idle_qq <= #TCQ 1'b1;
            pipe_tx_powerdown_qq <= #TCQ 2'b10;

        end 
        else 
        begin

            pipe_rx_char_is_k_q <= #TCQ pipe_rx_char_is_k_i;
            pipe_rx_data_q <= #TCQ pipe_rx_data_i;
            pipe_rx_valid_q <= #TCQ pipe_rx_valid_i;
            pipe_rx_chanisaligned_q <= #TCQ pipe_rx_chanisaligned_i;
            pipe_rx_status_q <= #TCQ pipe_rx_status_i;
            pipe_rx_phy_status_q <= #TCQ pipe_rx_phy_status_i;
            pipe_rx_elec_idle_q <= #TCQ pipe_rx_elec_idle_i;

            pipe_rx_polarity_q <= #TCQ pipe_rx_polarity_i;
            pipe_tx_compliance_q <= #TCQ pipe_tx_compliance_i;
            pipe_tx_char_is_k_q <= #TCQ pipe_tx_char_is_k_i;
            pipe_tx_data_q <= #TCQ pipe_tx_data_i;
            pipe_tx_elec_idle_q <= #TCQ pipe_tx_elec_idle_i;
            pipe_tx_powerdown_q <= #TCQ pipe_tx_powerdown_i;

            pipe_rx_char_is_k_qq <= #TCQ pipe_rx_char_is_k_q;
            pipe_rx_data_qq <= #TCQ pipe_rx_data_q;
            pipe_rx_valid_qq <= #TCQ pipe_rx_valid_q;
            pipe_rx_chanisaligned_qq <= #TCQ pipe_rx_chanisaligned_q;
            pipe_rx_status_qq <= #TCQ pipe_rx_status_q;
            pipe_rx_phy_status_qq <= #TCQ pipe_rx_phy_status_q;
            pipe_rx_elec_idle_qq <= #TCQ pipe_rx_elec_idle_q;

            pipe_rx_polarity_qq <= #TCQ pipe_rx_polarity_q;
            pipe_tx_compliance_qq <= #TCQ pipe_tx_compliance_q;
            pipe_tx_char_is_k_qq <= #TCQ pipe_tx_char_is_k_q;
            pipe_tx_data_qq <= #TCQ pipe_tx_data_q;
            pipe_tx_elec_idle_qq <= #TCQ pipe_tx_elec_idle_q;
            pipe_tx_powerdown_qq <= #TCQ pipe_tx_powerdown_q;

          end

        end

        assign pipe_rx_char_is_k_o = pipe_rx_char_is_k_qq;
        assign pipe_rx_data_o = pipe_rx_data_qq;
        assign pipe_rx_valid_o = pipe_rx_valid_qq;
        assign pipe_rx_chanisaligned_o = pipe_rx_chanisaligned_qq;
        assign pipe_rx_status_o = pipe_rx_status_qq;
        assign pipe_rx_phy_status_o = pipe_rx_phy_status_qq;
        assign pipe_rx_elec_idle_o = pipe_rx_elec_idle_qq;

        assign pipe_rx_polarity_o = pipe_rx_polarity_qq;
        assign pipe_tx_compliance_o = pipe_tx_compliance_qq;
        assign pipe_tx_char_is_k_o = pipe_tx_char_is_k_qq;
        assign pipe_tx_data_o = pipe_tx_data_qq;
        assign pipe_tx_elec_idle_o = pipe_tx_elec_idle_qq;
        assign pipe_tx_powerdown_o = pipe_tx_powerdown_qq;

    end // if (PIPE_PIPELINE_STAGES == 2)

    endgenerate

endmodule



`timescale 1ns/1ps
module model_ap2_tst_gt_top #
(
   parameter               LINK_CAP_MAX_LINK_WIDTH = 8,          // 1 - x1 , 2 - x2 , 4 - x4 , 8 - x8
   parameter               REF_CLK_FREQ            = 0,          // 0 - 100 MHz , 1 - 125 MHz , 2 - 250 MHz
   parameter               USER_CLK2_DIV2          = "FALSE",    // "FALSE" => user_clk2 = user_clk
                                                                 // "TRUE" => user_clk2 = user_clk/2, where user_clk = 500 or 250 MHz.
   parameter  integer      USER_CLK_FREQ           = 3,          // 0 - 31.25 MHz , 1 - 62.5 MHz , 2 - 125 MHz , 3 - 250 MHz , 4 - 500Mhz
   parameter               PL_FAST_TRAIN           = "FALSE",    // Simulation Speedup
   parameter               PCIE_EXT_CLK            = "FALSE",    // Use External Clocking
   parameter               PCIE_USE_MODE           = "1.0",      // 1.0 = K325T IES, 1.1 = VX485T IES, 3.0 = K325T GES
   parameter               PCIE_GT_DEVICE          = "GTX",      // Select the GT to use (GTP for Artix-7, GTX for K7/V7)
   parameter               PCIE_PLL_SEL            = "CPLL",     // Select the PLL (CPLL or QPLL)
   parameter               PCIE_ASYNC_EN           = "FALSE",    // Asynchronous Clocking Enable
   parameter               PCIE_TXBUF_EN           = "FALSE",    // Use the Tansmit Buffer
   parameter               PCIE_EXT_GT_COMMON      = "FALSE", 
   parameter               EXT_CH_GT_DRP           = "FALSE",  
   parameter               TX_MARGIN_FULL_0        = 7'b1001111, // 1000 mV
   parameter               TX_MARGIN_FULL_1        = 7'b1001110, // 950 mV
   parameter               TX_MARGIN_FULL_2        = 7'b1001101, // 900 mV
   parameter               TX_MARGIN_FULL_3        = 7'b1001100, // 850 mV
   parameter               TX_MARGIN_FULL_4        = 7'b1000011, // 400 mV
   parameter               TX_MARGIN_LOW_0         = 7'b1000101, // 500 mV
   parameter               TX_MARGIN_LOW_1         = 7'b1000110, // 450 mV
   parameter               TX_MARGIN_LOW_2         = 7'b1000011, // 400 mV
   parameter               TX_MARGIN_LOW_3         = 7'b1000010, // 350 mV
   parameter               TX_MARGIN_LOW_4         = 7'b1000000,   

   parameter               PCIE_CHAN_BOND          = 0,
   parameter               TCQ                     = 1           //synthesis warning solved: parameter declaration becomes local
)
(
   //-----------------------------------------------------------------------------------------------------------------//
   // pl ltssm
   input   wire [5:0]                pl_ltssm_state         ,
   // Pipe Per-Link Signals
   input   wire                      pipe_tx_rcvr_det       ,
   input   wire                      pipe_tx_reset          ,
   input   wire                      pipe_tx_rate           ,
   input   wire                      pipe_tx_deemph         ,
   input   wire [2:0]                pipe_tx_margin         ,
   input   wire                      pipe_tx_swing          ,

   //-----------------------------------------------------------------------------------------------------------------//
   // Pipe Per-Lane Signals                                                                                           //
   //-----------------------------------------------------------------------------------------------------------------//


   // Pipe Per-Lane Signals - Lane 0
   output  wire [ 1:0]               pipe_rx0_char_is_k     ,
   output  wire [15:0]               pipe_rx0_data          ,
   output  wire                      pipe_rx0_valid         ,
   output  wire                      pipe_rx0_chanisaligned ,
   output  wire [ 2:0]               pipe_rx0_status        ,
   output  wire                      pipe_rx0_phy_status    ,
   output  wire                      pipe_rx0_elec_idle     ,
   input   wire                      pipe_rx0_polarity      ,
   input   wire                      pipe_tx0_compliance    ,
   input   wire [ 1:0]               pipe_tx0_char_is_k     ,
   input   wire [15:0]               pipe_tx0_data          ,
   input   wire                      pipe_tx0_elec_idle     ,
   input   wire [ 1:0]               pipe_tx0_powerdown     ,

   // Pipe Per-Lane Signals - Lane 1
   output  wire [ 1:0]               pipe_rx1_char_is_k     ,
   output  wire [15:0]               pipe_rx1_data          ,
   output  wire                      pipe_rx1_valid         ,
   output  wire                      pipe_rx1_chanisaligned ,
   output  wire [ 2:0]               pipe_rx1_status        ,
   output  wire                      pipe_rx1_phy_status    ,
   output  wire                      pipe_rx1_elec_idle     ,
   input   wire                      pipe_rx1_polarity      ,
   input   wire                      pipe_tx1_compliance    ,
   input   wire [ 1:0]               pipe_tx1_char_is_k     ,
   input   wire [15:0]               pipe_tx1_data          ,
   input   wire                      pipe_tx1_elec_idle     ,
   input   wire [ 1:0]               pipe_tx1_powerdown     ,

   // Pipe Per-Lane Signals - Lane 2
   output  wire [ 1:0]               pipe_rx2_char_is_k     ,
   output  wire [15:0]               pipe_rx2_data          ,
   output  wire                      pipe_rx2_valid         ,
   output  wire                      pipe_rx2_chanisaligned ,
   output  wire [ 2:0]               pipe_rx2_status        ,
   output  wire                      pipe_rx2_phy_status    ,
   output  wire                      pipe_rx2_elec_idle     ,
   input   wire                      pipe_rx2_polarity      ,
   input   wire                      pipe_tx2_compliance    ,
   input   wire [ 1:0]               pipe_tx2_char_is_k     ,
   input   wire [15:0]               pipe_tx2_data          ,
   input   wire                      pipe_tx2_elec_idle     ,
   input   wire [ 1:0]               pipe_tx2_powerdown     ,

   // Pipe Per-Lane Signals - Lane 3
   output  wire [ 1:0]               pipe_rx3_char_is_k     ,
   output  wire [15:0]               pipe_rx3_data          ,
   output  wire                      pipe_rx3_valid         ,
   output  wire                      pipe_rx3_chanisaligned ,
   output  wire [ 2:0]               pipe_rx3_status        ,
   output  wire                      pipe_rx3_phy_status    ,
   output  wire                      pipe_rx3_elec_idle     ,
   input   wire                      pipe_rx3_polarity      ,
   input   wire                      pipe_tx3_compliance    ,
   input   wire [ 1:0]               pipe_tx3_char_is_k     ,
   input   wire [15:0]               pipe_tx3_data          ,
   input   wire                      pipe_tx3_elec_idle     ,
   input   wire [ 1:0]               pipe_tx3_powerdown     ,

   // Pipe Per-Lane Signals - Lane 4
   output  wire [ 1:0]               pipe_rx4_char_is_k     ,
   output  wire [15:0]               pipe_rx4_data          ,
   output  wire                      pipe_rx4_valid         ,
   output  wire                      pipe_rx4_chanisaligned ,
   output  wire [ 2:0]               pipe_rx4_status        ,
   output  wire                      pipe_rx4_phy_status    ,
   output  wire                      pipe_rx4_elec_idle     ,
   input   wire                      pipe_rx4_polarity      ,
   input   wire                      pipe_tx4_compliance    ,
   input   wire [ 1:0]               pipe_tx4_char_is_k     ,
   input   wire [15:0]               pipe_tx4_data          ,
   input   wire                      pipe_tx4_elec_idle     ,
   input   wire [ 1:0]               pipe_tx4_powerdown     ,

   // Pipe Per-Lane Signals - Lane 5
   output  wire [ 1:0]               pipe_rx5_char_is_k     ,
   output  wire [15:0]               pipe_rx5_data          ,
   output  wire                      pipe_rx5_valid         ,
   output  wire                      pipe_rx5_chanisaligned ,
   output  wire [ 2:0]               pipe_rx5_status        ,
   output  wire                      pipe_rx5_phy_status    ,
   output  wire                      pipe_rx5_elec_idle     ,
   input   wire                      pipe_rx5_polarity      ,
   input   wire                      pipe_tx5_compliance    ,
   input   wire [ 1:0]               pipe_tx5_char_is_k     ,
   input   wire [15:0]               pipe_tx5_data          ,
   input   wire                      pipe_tx5_elec_idle     ,
   input   wire [ 1:0]               pipe_tx5_powerdown     ,

   // Pipe Per-Lane Signals - Lane 6
   output  wire [ 1:0]               pipe_rx6_char_is_k     ,
   output  wire [15:0]               pipe_rx6_data          ,
   output  wire                      pipe_rx6_valid         ,
   output  wire                      pipe_rx6_chanisaligned ,
   output  wire [ 2:0]               pipe_rx6_status        ,
   output  wire                      pipe_rx6_phy_status    ,
   output  wire                      pipe_rx6_elec_idle     ,
   input   wire                      pipe_rx6_polarity      ,
   input   wire                      pipe_tx6_compliance    ,
   input   wire [ 1:0]               pipe_tx6_char_is_k     ,
   input   wire [15:0]               pipe_tx6_data          ,
   input   wire                      pipe_tx6_elec_idle     ,
   input   wire [ 1:0]               pipe_tx6_powerdown     ,

   // Pipe Per-Lane Signals - Lane 7
   output  wire [ 1:0]               pipe_rx7_char_is_k     ,
   output  wire [15:0]               pipe_rx7_data          ,
   output  wire                      pipe_rx7_valid         ,
   output  wire                      pipe_rx7_chanisaligned ,
   output  wire [ 2:0]               pipe_rx7_status        ,
   output  wire                      pipe_rx7_phy_status    ,
   output  wire                      pipe_rx7_elec_idle     ,
   input   wire                      pipe_rx7_polarity      ,
   input   wire                      pipe_tx7_compliance    ,
   input   wire [ 1:0]               pipe_tx7_char_is_k     ,
   input   wire [15:0]               pipe_tx7_data          ,
   input   wire                      pipe_tx7_elec_idle     ,
   input   wire [ 1:0]               pipe_tx7_powerdown     ,

   // PCI Express signals
   output  wire [ (LINK_CAP_MAX_LINK_WIDTH-1):0] pci_exp_txn            ,
   output  wire [ (LINK_CAP_MAX_LINK_WIDTH-1):0] pci_exp_txp            ,
   input   wire [ (LINK_CAP_MAX_LINK_WIDTH-1):0] pci_exp_rxn            ,
   input   wire [ (LINK_CAP_MAX_LINK_WIDTH-1):0] pci_exp_rxp            ,

   // Non PIPE signals
   input   wire                                  sys_clk                ,
   input   wire                                  sys_rst_n              ,
   input   wire                                  PIPE_MMCM_RST_N        ,
   output  wire                                  pipe_clk               ,
   output  wire                                  user_clk               ,
   output  wire                                  user_clk2              ,

//----------- Shared Logic Internal--------------------------------------

  output                                        INT_PCLK_OUT_SLAVE,     // PCLK       | PCLK
  output                                        INT_RXUSRCLK_OUT,       // RXUSERCLK
  output  [(LINK_CAP_MAX_LINK_WIDTH-1):0]       INT_RXOUTCLK_OUT,       // RX recovered clock
  output                                        INT_DCLK_OUT,           // DCLK       | DCLK
  output                                        INT_USERCLK1_OUT,       // Optional user clock
  output                                        INT_USERCLK2_OUT,       // Optional user clock
  output                                        INT_OOBCLK_OUT,         // OOB        | OOB
  output                                        INT_MMCM_LOCK_OUT,      // Async      | Async
  output  [1:0]                                 INT_QPLLLOCK_OUT,
  output  [1:0]                                 INT_QPLLOUTCLK_OUT,
  output  [1:0]                                 INT_QPLLOUTREFCLK_OUT,
  input   [(LINK_CAP_MAX_LINK_WIDTH-1):0]       INT_PCLK_SEL_SLAVE,

  // Shared Logic External

 //---------- External GT COMMON Ports ----------------------
  input   [11:0]                                qpll_drp_crscode,
  input   [17:0]                                qpll_drp_fsm,
  input   [1:0]                                 qpll_drp_done,
  input   [1:0]                                 qpll_drp_reset,
  input   [1:0]                                 qpll_qplllock,
  input   [1:0]                                 qpll_qplloutclk,
  input   [1:0]                                 qpll_qplloutrefclk,
  output                                        qpll_qplld,
  output  [1:0]                                 qpll_qpllreset,
  output                                        qpll_drp_clk,
  output                                        qpll_drp_rst_n,
  output                                        qpll_drp_ovrd,
  output                                        qpll_drp_gen3,
  output                                        qpll_drp_start,

  //---------- External Clock Ports ----------------------
  input                                         PIPE_PCLK_IN,           // PCLK       | PCLK
  input                                         PIPE_RXUSRCLK_IN,       // RXUSERCLK
  input  [LINK_CAP_MAX_LINK_WIDTH-1:0]          PIPE_RXOUTCLK_IN,       // RX recovered clock
  input                                         PIPE_DCLK_IN,           // DCLK       | DCLK
  input                                         PIPE_USERCLK1_IN,       // Optional user clock
  input                                         PIPE_USERCLK2_IN,       // Optional user clock
  input                                         PIPE_OOBCLK_IN,         // OOB        | OOB
  input                                         PIPE_MMCM_LOCK_IN,      // Async      | Async
  output                                        PIPE_TXOUTCLK_OUT,      // PCLK       | PCLK
  output [LINK_CAP_MAX_LINK_WIDTH-1:0]          PIPE_RXOUTCLK_OUT,      // RX recovered clock (for debug only)
  output [LINK_CAP_MAX_LINK_WIDTH-1:0]          PIPE_PCLK_SEL_OUT,      // PCLK       | PCLK
  output                                        PIPE_GEN3_OUT ,          // PCLK       | PCLK

//-----------TRANSCEIVER DEBUG--------------------------------

  output      [4:0]                             PIPE_RST_FSM,
  output      [11:0]                            PIPE_QRST_FSM,
  output      [(LINK_CAP_MAX_LINK_WIDTH*5)-1:0] PIPE_RATE_FSM,
  output      [(LINK_CAP_MAX_LINK_WIDTH*6)-1:0] PIPE_SYNC_FSM_TX,
  output      [(LINK_CAP_MAX_LINK_WIDTH*7)-1:0] PIPE_SYNC_FSM_RX,
  output      [(LINK_CAP_MAX_LINK_WIDTH*7)-1:0] PIPE_DRP_FSM,

  output                                        PIPE_RST_IDLE,
  output                                        PIPE_QRST_IDLE,
  output                                        PIPE_RATE_IDLE,
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_EYESCANDATAERROR,
  output     [(LINK_CAP_MAX_LINK_WIDTH*3)-1:0]  PIPE_RXSTATUS,
  output     [(LINK_CAP_MAX_LINK_WIDTH*15)-1:0] PIPE_DMONITOROUT,

  //---------- Debug Ports -------------------------------
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_CPLL_LOCK,
  output     [(LINK_CAP_MAX_LINK_WIDTH-1)>>2:0] PIPE_QPLL_LOCK,
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_RXPMARESETDONE,       
  output     [(LINK_CAP_MAX_LINK_WIDTH*3)-1:0]  PIPE_RXBUFSTATUS,         
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_TXPHALIGNDONE,       
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_TXPHINITDONE,        
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_TXDLYSRESETDONE,    
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_RXPHALIGNDONE,      
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_RXDLYSRESETDONE,     
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_RXSYNCDONE,       
  output     [(LINK_CAP_MAX_LINK_WIDTH*8)-1:0]  PIPE_RXDISPERR,       
  output     [(LINK_CAP_MAX_LINK_WIDTH*8)-1:0]  PIPE_RXNOTINTABLE,      
  output     [(LINK_CAP_MAX_LINK_WIDTH)-1:0]    PIPE_RXCOMMADET,        

  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_0,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_1,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_2,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_3,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_4,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_5,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_6,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_7,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_8,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_DEBUG_9,
  output      [31:0]                            PIPE_DEBUG,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_JTAG_RDY,

  input       [ 2:0]                            PIPE_TXPRBSSEL,
  input       [ 2:0]                            PIPE_RXPRBSSEL,
  input                                         PIPE_TXPRBSFORCEERR,
  input                                         PIPE_RXPRBSCNTRESET,
  input       [ 2:0]                            PIPE_LOOPBACK,
  output      [LINK_CAP_MAX_LINK_WIDTH-1:0]     PIPE_RXPRBSERR,

  //-----------Channel DRP----------------------------------------
  output                                          ext_ch_gt_drpclk,
  input        [(LINK_CAP_MAX_LINK_WIDTH*9)-1:0] ext_ch_gt_drpaddr,
  input        [LINK_CAP_MAX_LINK_WIDTH-1:0]     ext_ch_gt_drpen,
  input        [(LINK_CAP_MAX_LINK_WIDTH*16)-1:0]ext_ch_gt_drpdi,
  input        [LINK_CAP_MAX_LINK_WIDTH-1:0]     ext_ch_gt_drpwe,

  output       [(LINK_CAP_MAX_LINK_WIDTH*16)-1:0]ext_ch_gt_drpdo,
  output       [LINK_CAP_MAX_LINK_WIDTH-1:0]     ext_ch_gt_drprdy,

  output  wire                      phy_rdy_n
);


  localparam                         USERCLK2_FREQ   =  (USER_CLK2_DIV2 == "FALSE") ? USER_CLK_FREQ :
                                                        (USER_CLK_FREQ == 4) ? 3 :
                                                        (USER_CLK_FREQ == 3) ? 2 :
                                                         USER_CLK_FREQ;

  localparam                         PCIE_LPM_DFE    = (PL_FAST_TRAIN == "TRUE") ? "DFE" : "LPM";
  localparam                         PCIE_LINK_SPEED = (PL_FAST_TRAIN == "TRUE") ? 2 : 3;

  // The parameter PCIE_OOBCLK_MODE_ENABLE value should be "0" for simulation and for synthesis it should be 1
  //localparam                         PCIE_OOBCLK_MODE_ENABLE = (PL_FAST_TRAIN == "TRUE") ? 0 : 1;  
  localparam                         PCIE_OOBCLK_MODE_ENABLE = 1;  

  localparam              PCIE_TX_EIDLE_ASSERT_DELAY = (PL_FAST_TRAIN == "TRUE") ? 3'd4 : 3'd2;

  wire [  7:0]                       gt_rx_phy_status_wire        ;
  wire [  7:0]                       gt_rxchanisaligned_wire      ;
  wire [ 31:0]                       gt_rx_data_k_wire            ;
  wire [255:0]                       gt_rx_data_wire              ;
  wire [  7:0]                       gt_rx_elec_idle_wire         ;
  wire [ 23:0]                       gt_rx_status_wire            ;
  wire [  7:0]                       gt_rx_valid_wire             ;
  wire [  7:0]                       gt_rx_polarity               ;
  wire [ 15:0]                       gt_power_down                ;
  wire [  7:0]                       gt_tx_char_disp_mode         ;
  wire [ 31:0]                       gt_tx_data_k                 ;
  wire [255:0]                       gt_tx_data                   ;
  wire                               gt_tx_detect_rx_loopback     ;
  wire [  7:0]                       gt_tx_elec_idle              ;
  wire [  7:0]                       gt_rx_elec_idle_reset        ;
  wire [LINK_CAP_MAX_LINK_WIDTH-1:0] phystatus_rst                ;
  wire                               clock_locked                 ;

  wire [  7:0]                       gt_rx_phy_status_wire_filter ;
  wire [ 31:0]                       gt_rx_data_k_wire_filter     ;
  wire [255:0]                       gt_rx_data_wire_filter       ;
  wire [  7:0]                       gt_rx_elec_idle_wire_filter  ;
  wire [ 23:0]                       gt_rx_status_wire_filter     ;
  wire [  7:0]                       gt_rx_valid_wire_filter      ;

  wire [LINK_CAP_MAX_LINK_WIDTH-1:0] gt_eyescandataerror          ;
  wire                               pipe_clk_int;
  reg                                phy_rdy_n_int;

  reg                                reg_clock_locked;
  wire                               all_phystatus_rst;

reg [5:0] pl_ltssm_state_q;

always @(posedge pipe_clk_int or negedge clock_locked) begin

  if (!clock_locked)
    pl_ltssm_state_q <= #TCQ 6'b0;
  else
    pl_ltssm_state_q <= #TCQ pl_ltssm_state;

end

  assign pipe_clk = pipe_clk_int ;

  wire                               plm_in_l0 = (pl_ltssm_state_q == 6'h16);
  wire                               plm_in_rl = (pl_ltssm_state_q == 6'h1c);
  wire                               plm_in_dt = (pl_ltssm_state_q == 6'h2d);
  wire                               plm_in_rs = (pl_ltssm_state_q == 6'h1f);

//-------------RX FILTER Instantiation----------------------------------------------------------//
genvar i;
generate for (i=0; i<LINK_CAP_MAX_LINK_WIDTH; i=i+1)
 begin : gt_rx_valid_filter

model_ap2_tst_gt_rx_valid_filter_7x # (
     .CLK_COR_MIN_LAT(28)
   )
   model_ap2_tst_GT_RX_VALID_FILTER_7x_inst (

     .USER_RXCHARISK   ( gt_rx_data_k_wire [(2*i)+1 + (2*i):(2*i)+ (2*i)] ),           //O
     .USER_RXDATA      ( gt_rx_data_wire [(16*i)+15+(16*i) :(16*i)+0 + (16*i)] ),      //O
     .USER_RXVALID     ( gt_rx_valid_wire [i] ),                                       //O
     .USER_RXELECIDLE  ( gt_rx_elec_idle_wire [i] ),                                   //O
     .USER_RX_STATUS   ( gt_rx_status_wire [(3*i)+2:(3*i)] ),                          //O
     .USER_RX_PHY_STATUS ( gt_rx_phy_status_wire [i] ),                                //O

     .GT_RXCHARISK     ( gt_rx_data_k_wire_filter [(2*i)+1+ (2*i):2*i+ (2*i)] ),       //I
     .GT_RXDATA        ( gt_rx_data_wire_filter [(16*i)+15+(16*i) :(16*i)+0+(16*i)] ), //I
     .GT_RXVALID       ( gt_rx_valid_wire_filter [i] ),                                //I
     .GT_RXELECIDLE    ( gt_rx_elec_idle_wire_filter [i] ),                            //I
     .GT_RX_STATUS     ( gt_rx_status_wire_filter [(3*i)+2:(3*i)] ),                   //I
     .GT_RX_PHY_STATUS ( gt_rx_phy_status_wire_filter [i] ),

     .PLM_IN_L0        ( plm_in_l0 ),                                                  //I
     .PLM_IN_RS        ( plm_in_rs ),                                                  //I
     .USER_CLK         ( pipe_clk_int ),                                               //I
     .RESET            ( phy_rdy_n_int )                                               //I
   );


 end
endgenerate

  //---------- GT Instantiation ---------------------------------------------------------------
model_ap2_tst_pipe_wrapper #
  (
    .PCIE_SIM_MODE                  ( PL_FAST_TRAIN ),
 
    // synthesis translate_off
    .PCIE_SIM_SPEEDUP               ( "TRUE" ),
    // synthesis translate_on

    .PCIE_EXT_CLK                   ( PCIE_EXT_CLK ),
    .PCIE_TXBUF_EN                  ( PCIE_TXBUF_EN ),
    .PCIE_EXT_GT_COMMON             ( PCIE_EXT_GT_COMMON ),
    .EXT_CH_GT_DRP                  ( EXT_CH_GT_DRP ),
    .TX_MARGIN_FULL_0               (TX_MARGIN_FULL_0),                          
    .TX_MARGIN_FULL_1               (TX_MARGIN_FULL_1),                          
    .TX_MARGIN_FULL_2               (TX_MARGIN_FULL_2),                          
    .TX_MARGIN_FULL_3               (TX_MARGIN_FULL_3),                          
    .TX_MARGIN_FULL_4               (TX_MARGIN_FULL_4),                          
    .TX_MARGIN_LOW_0                (TX_MARGIN_LOW_0),                          
    .TX_MARGIN_LOW_1                (TX_MARGIN_LOW_1),                          
    .TX_MARGIN_LOW_2                (TX_MARGIN_LOW_2),                          
    .TX_MARGIN_LOW_3                (TX_MARGIN_LOW_3),                          
    .TX_MARGIN_LOW_4                (TX_MARGIN_LOW_4),
    .PCIE_ASYNC_EN                  ( PCIE_ASYNC_EN ),
    .PCIE_CHAN_BOND                 ( PCIE_CHAN_BOND ),
    .PCIE_PLL_SEL                   ( PCIE_PLL_SEL ),
    .PCIE_GT_DEVICE                 ( PCIE_GT_DEVICE ),
    .PCIE_USE_MODE                  ( PCIE_USE_MODE ),
    .PCIE_LANE                      ( LINK_CAP_MAX_LINK_WIDTH ),
    .PCIE_LPM_DFE                   ( PCIE_LPM_DFE ),
    .PCIE_LINK_SPEED                ( PCIE_LINK_SPEED ),
    .PCIE_TX_EIDLE_ASSERT_DELAY     ( PCIE_TX_EIDLE_ASSERT_DELAY ),
    .PCIE_OOBCLK_MODE               ( PCIE_OOBCLK_MODE_ENABLE ),
    .PCIE_REFCLK_FREQ               ( REF_CLK_FREQ ),
    .PCIE_USERCLK1_FREQ             ( USER_CLK_FREQ +1 ),
    .PCIE_USERCLK2_FREQ             ( USERCLK2_FREQ +1 )

  ) model_ap2_tst_pipe_wrapper_i (

    //---------- PIPE Clock & Reset Ports ------------------
    .PIPE_CLK                        ( sys_clk ),
    .PIPE_RESET_N                    ( sys_rst_n ),
    .PIPE_PCLK                       ( pipe_clk_int ),

    //---------- PIPE TX Data Ports ------------------
    .PIPE_TXDATA                    ( gt_tx_data[((32*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_TXDATAK                   ( gt_tx_data_k[((4*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),

    .PIPE_TXP                       ( pci_exp_txp[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_TXN                       ( pci_exp_txn[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),

    //---------- PIPE RX Data Ports ------------------
    .PIPE_RXP                       ( pci_exp_rxp[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_RXN                       ( pci_exp_rxn[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),

    .PIPE_RXDATA                    ( gt_rx_data_wire_filter[((32*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_RXDATAK                   ( gt_rx_data_k_wire_filter[((4*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),

    //---------- PIPE Command Ports ------------------
    .PIPE_TXDETECTRX                ( gt_tx_detect_rx_loopback ),
    .PIPE_TXELECIDLE                ( gt_tx_elec_idle[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_TXCOMPLIANCE              ( gt_tx_char_disp_mode[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_RXPOLARITY                ( gt_rx_polarity[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_POWERDOWN                 ( gt_power_down[((2*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_RATE                      ( {1'b0,pipe_tx_rate} ),

    //---------- PIPE Electrical Command Ports ------------------
    .PIPE_TXMARGIN                  ( pipe_tx_margin[2:0] ),
    .PIPE_TXSWING                   ( pipe_tx_swing ),
    .PIPE_TXDEEMPH                  ( {(LINK_CAP_MAX_LINK_WIDTH){pipe_tx_deemph}}),
    .PIPE_TXEQ_CONTROL              ( {2*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_TXEQ_PRESET               ( {4*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_TXEQ_PRESET_DEFAULT       ( {4*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),

    .PIPE_RXEQ_CONTROL              ( {2*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_PRESET               ( {3*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_LFFS                 ( {6*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_TXPRESET             ( {4*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_USER_EN              ( {1*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_USER_TXCOEFF         ( {18*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_RXEQ_USER_MODE            ( {1*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_TXEQ_COEFF                ( ),
    .PIPE_TXEQ_DEEMPH               ( {6*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),
    .PIPE_TXEQ_FS                   ( ),
    .PIPE_TXEQ_LF                   ( ),
    .PIPE_TXEQ_DONE                 ( ),

    .PIPE_RXEQ_NEW_TXCOEFF          ( ),
    .PIPE_RXEQ_LFFS_SEL             ( ),
    .PIPE_RXEQ_ADAPT_DONE           ( ),
    .PIPE_RXEQ_DONE                 ( ),

    //---------- PIPE Status Ports -------------------
    .PIPE_RXVALID                   ( gt_rx_valid_wire_filter[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_PHYSTATUS                 ( gt_rx_phy_status_wire_filter[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_PHYSTATUS_RST             ( phystatus_rst ),
    .PIPE_RXELECIDLE                ( gt_rx_elec_idle_wire_filter[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_EYESCANDATAERROR          ( gt_eyescandataerror[((LINK_CAP_MAX_LINK_WIDTH)-1):0] ),
    .PIPE_RXSTATUS                  ( gt_rx_status_wire_filter[((3*LINK_CAP_MAX_LINK_WIDTH)-1):0] ),

    .INT_PCLK_OUT_SLAVE             (INT_PCLK_OUT_SLAVE   ),           
    .INT_RXUSRCLK_OUT               (INT_RXUSRCLK_OUT     ),    
    .INT_RXOUTCLK_OUT               (INT_RXOUTCLK_OUT     ),         
    .INT_DCLK_OUT                   (INT_DCLK_OUT         ),           
    .INT_USERCLK1_OUT               (INT_USERCLK1_OUT     ),      
    .INT_USERCLK2_OUT               (INT_USERCLK2_OUT     ),       
    .INT_OOBCLK_OUT                 (INT_OOBCLK_OUT       ),     
    .INT_MMCM_LOCK_OUT              (INT_MMCM_LOCK_OUT    ),        
    .INT_QPLLLOCK_OUT               (INT_QPLLLOCK_OUT     ),        
    .INT_QPLLOUTCLK_OUT             (INT_QPLLOUTCLK_OUT   ),        
    .INT_QPLLOUTREFCLK_OUT          (INT_QPLLOUTREFCLK_OUT),         
    .INT_PCLK_SEL_SLAVE             (INT_PCLK_SEL_SLAVE   ),    
    //---------- PIPE User Ports ---------------------------
    .PIPE_MMCM_RST_N                ( PIPE_MMCM_RST_N ),        // Async      | Async

    .PIPE_RXSLIDE                   ( {1*LINK_CAP_MAX_LINK_WIDTH{1'b0}} ),

    .PIPE_PCLK_LOCK                 ( clock_locked ),
    .PIPE_RXCDRLOCK                 ( ),
    .PIPE_USERCLK1                  ( user_clk ),
    .PIPE_USERCLK2                  ( user_clk2 ),
    .PIPE_RXUSRCLK                  ( ),

    .PIPE_RXOUTCLK                  ( ),
    .PIPE_TXSYNC_DONE               ( ),
    .PIPE_RXSYNC_DONE               ( ),
    .PIPE_GEN3_RDY                  ( ),
    .PIPE_RXCHANISALIGNED           ( gt_rxchanisaligned_wire[LINK_CAP_MAX_LINK_WIDTH-1:0] ),
    .PIPE_ACTIVE_LANE               ( ),

    //---------- External Clock Ports ---------------------------
    .PIPE_PCLK_IN                   ( PIPE_PCLK_IN ),
    .PIPE_RXUSRCLK_IN               ( PIPE_RXUSRCLK_IN ),

    .PIPE_RXOUTCLK_IN               ( PIPE_RXOUTCLK_IN ),
    .PIPE_DCLK_IN                   ( PIPE_DCLK_IN ),
    .PIPE_USERCLK1_IN               ( PIPE_USERCLK1_IN ),
    .PIPE_USERCLK2_IN               ( PIPE_USERCLK2_IN ),
    .PIPE_OOBCLK_IN                 ( PIPE_OOBCLK_IN ),
    .PIPE_JTAG_EN                   ( 1'b0 ),
    .PIPE_JTAG_RDY                  ( PIPE_JTAG_RDY ),
    .PIPE_MMCM_LOCK_IN              ( PIPE_MMCM_LOCK_IN ),

    .PIPE_TXOUTCLK_OUT              ( PIPE_TXOUTCLK_OUT ),
    .PIPE_RXOUTCLK_OUT              ( PIPE_RXOUTCLK_OUT ),
    .PIPE_PCLK_SEL_OUT              ( PIPE_PCLK_SEL_OUT ),
    .PIPE_GEN3_OUT                  ( PIPE_GEN3_OUT ),
 //--------TRANSCEIVER DEBUG EOU------------------
   .EXT_CH_GT_DRPCLK          (ext_ch_gt_drpclk),
   .EXT_CH_GT_DRPADDR         (ext_ch_gt_drpaddr),
   .EXT_CH_GT_DRPEN           (ext_ch_gt_drpen),
   .EXT_CH_GT_DRPDI           (ext_ch_gt_drpdi),
   .EXT_CH_GT_DRPWE           (ext_ch_gt_drpwe),
   .EXT_CH_GT_DRPDO           (ext_ch_gt_drpdo),
   .EXT_CH_GT_DRPRDY          (ext_ch_gt_drprdy),

   //---------- External GT COMMON Ports ----------------------
    .QPLL_DRP_CRSCODE         ( qpll_drp_crscode ),
    .QPLL_DRP_FSM             ( qpll_drp_fsm ),
    .QPLL_DRP_DONE            ( qpll_drp_done ),
    .QPLL_DRP_RESET           ( qpll_drp_reset ),
    .QPLL_QPLLLOCK            ( qpll_qplllock ),
    .QPLL_QPLLOUTCLK          ( qpll_qplloutclk ),
    .QPLL_QPLLOUTREFCLK       ( qpll_qplloutrefclk ),
    .QPLL_QPLLPD              ( qpll_qplld ),
    .QPLL_QPLLRESET           ( qpll_qpllreset ),
    .QPLL_DRP_CLK             ( qpll_drp_clk ),
    .QPLL_DRP_RST_N           ( qpll_drp_rst_n ),
    .QPLL_DRP_OVRD            ( qpll_drp_ovrd ),
    .QPLL_DRP_GEN3            ( qpll_drp_gen3 ),
    .QPLL_DRP_START           ( qpll_drp_start ),

  //---------- TRANSCEIVER DEBUG -----------------------
    .PIPE_TXPRBSSEL           ( PIPE_TXPRBSSEL ),
    .PIPE_RXPRBSSEL           ( PIPE_RXPRBSSEL ),
    .PIPE_TXPRBSFORCEERR      ( PIPE_TXPRBSFORCEERR ),
    .PIPE_RXPRBSCNTRESET      ( PIPE_RXPRBSCNTRESET ),
    .PIPE_LOOPBACK            ( PIPE_LOOPBACK ),

    .PIPE_RXPRBSERR           ( PIPE_RXPRBSERR ),

    .PIPE_RST_FSM             ( PIPE_RST_FSM ),
    .PIPE_QRST_FSM            ( PIPE_QRST_FSM ),
    .PIPE_RATE_FSM            ( PIPE_RATE_FSM ),
    .PIPE_SYNC_FSM_TX         ( PIPE_SYNC_FSM_TX ),
    .PIPE_SYNC_FSM_RX         ( PIPE_SYNC_FSM_RX ),
    .PIPE_QDRP_FSM            ( ),
    .PIPE_RXEQ_FSM            ( ),
    .PIPE_TXEQ_FSM            ( ),
    .PIPE_DRP_FSM             ( PIPE_DRP_FSM ),

    .PIPE_RST_IDLE            ( PIPE_RST_IDLE ),
    .PIPE_QRST_IDLE           ( PIPE_QRST_IDLE ),
    .PIPE_RATE_IDLE           ( PIPE_RATE_IDLE ),

    .PIPE_CPLL_LOCK           ( PIPE_CPLL_LOCK ),
    .PIPE_QPLL_LOCK           ( PIPE_QPLL_LOCK ),
    .PIPE_RXPMARESETDONE      ( PIPE_RXPMARESETDONE ),       
    .PIPE_RXBUFSTATUS         ( PIPE_RXBUFSTATUS    ),         
    .PIPE_TXPHALIGNDONE       ( PIPE_TXPHALIGNDONE  ),       
    .PIPE_TXPHINITDONE        ( PIPE_TXPHINITDONE   ),        
    .PIPE_TXDLYSRESETDONE     ( PIPE_TXDLYSRESETDONE),    
    .PIPE_RXPHALIGNDONE       ( PIPE_RXPHALIGNDONE  ),      
    .PIPE_RXDLYSRESETDONE     ( PIPE_RXDLYSRESETDONE),     
    .PIPE_RXSYNCDONE          ( PIPE_RXSYNCDONE     ),       
    .PIPE_RXDISPERR           ( PIPE_RXDISPERR      ),       
    .PIPE_RXNOTINTABLE        ( PIPE_RXNOTINTABLE   ),      
    .PIPE_RXCOMMADET          ( PIPE_RXCOMMADET     ),        
    //---------- Debug Ports -------------------------------
    .PIPE_DEBUG_0             ( PIPE_DEBUG_0  ),
    .PIPE_DEBUG_1             ( PIPE_DEBUG_1  ),
    .PIPE_DEBUG_2             ( PIPE_DEBUG_2  ),
    .PIPE_DEBUG_3             ( PIPE_DEBUG_3  ),
    .PIPE_DEBUG_4             ( PIPE_DEBUG_4  ),
    .PIPE_DEBUG_5             ( PIPE_DEBUG_5  ),
    .PIPE_DEBUG_6             ( PIPE_DEBUG_6  ),
    .PIPE_DEBUG_7             ( PIPE_DEBUG_7  ),
    .PIPE_DEBUG_8             ( PIPE_DEBUG_8  ),
    .PIPE_DEBUG_9             ( PIPE_DEBUG_9  ),
    .PIPE_DEBUG               ( PIPE_DEBUG    ),
    .PIPE_DMONITOROUT         ( PIPE_DMONITOROUT )
);

assign PIPE_RXSTATUS = gt_rx_status_wire_filter;
assign PIPE_EYESCANDATAERROR = gt_eyescandataerror;

assign pipe_rx0_phy_status = gt_rx_phy_status_wire[0] ;
assign pipe_rx1_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 2 ) ? gt_rx_phy_status_wire[1] : 1'b0;
assign pipe_rx2_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_phy_status_wire[2] : 1'b0;
assign pipe_rx3_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_phy_status_wire[3] : 1'b0;
assign pipe_rx4_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_phy_status_wire[4] : 1'b0;
assign pipe_rx5_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_phy_status_wire[5] : 1'b0;
assign pipe_rx6_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_phy_status_wire[6] : 1'b0;
assign pipe_rx7_phy_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_phy_status_wire[7] : 1'b0;

assign pipe_rx0_chanisaligned = gt_rxchanisaligned_wire[0];
assign pipe_rx1_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 2 ) ? gt_rxchanisaligned_wire[1] : 1'b0 ;
assign pipe_rx2_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rxchanisaligned_wire[2] : 1'b0 ;
assign pipe_rx3_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rxchanisaligned_wire[3] : 1'b0 ;
assign pipe_rx4_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rxchanisaligned_wire[4] : 1'b0 ;
assign pipe_rx5_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rxchanisaligned_wire[5] : 1'b0 ;
assign pipe_rx6_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rxchanisaligned_wire[6] : 1'b0 ;
assign pipe_rx7_chanisaligned = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rxchanisaligned_wire[7] : 1'b0 ;

//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<
//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<

generate
  if (LINK_CAP_MAX_LINK_WIDTH == 1)
   begin : rx_link_width_x1

     assign pipe_rx0_char_is_k =  {gt_rx_data_k_wire[1], gt_rx_data_k_wire[0]};
     assign pipe_rx1_char_is_k =  2'b0 ;
     assign pipe_rx2_char_is_k =  2'b0 ;
     assign pipe_rx3_char_is_k =  2'b0 ;
     assign pipe_rx4_char_is_k =  2'b0 ;
     assign pipe_rx5_char_is_k =  2'b0 ;
     assign pipe_rx6_char_is_k =  2'b0 ;
     assign pipe_rx7_char_is_k =  2'b0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_k_wire[3:2]   = 2'b0; 
     assign gt_rx_data_k_wire[5:4]   = 2'b0; 
     assign gt_rx_data_k_wire[7:6]   = 2'b0; 
     assign gt_rx_data_k_wire[9:8]   = 2'b0; 
     assign gt_rx_data_k_wire[11:10] = 2'b0; 
     assign gt_rx_data_k_wire[13:12] = 2'b0; 
     assign gt_rx_data_k_wire[15:14] = 2'b0; 
     assign gt_rx_data_k_wire[17:16] = 2'b0; 
     assign gt_rx_data_k_wire[19:18] = 2'b0; 
     assign gt_rx_data_k_wire[21:20] = 2'b0; 
     assign gt_rx_data_k_wire[23:22] = 2'b0; 
     assign gt_rx_data_k_wire[25:24] = 2'b0; 
     assign gt_rx_data_k_wire[27:26] = 2'b0; 
     assign gt_rx_data_k_wire[29:28] = 2'b0; 
     assign gt_rx_data_k_wire[31:30] = 2'b0; 

     assign pipe_rx0_data = {gt_rx_data_wire[ 15: 8], gt_rx_data_wire[ 7: 0]};
     assign pipe_rx1_data = 16'h0 ;
     assign pipe_rx2_data = 16'h0 ;
     assign pipe_rx3_data = 16'h0 ;
     assign pipe_rx4_data = 16'h0 ;
     assign pipe_rx5_data = 16'h0 ;
     assign pipe_rx6_data = 16'h0 ;
     assign pipe_rx7_data = 16'h0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_wire[31:16]   = 16'b0; 
     assign gt_rx_data_wire[47:32]   = 16'b0; 
     assign gt_rx_data_wire[63:48]   = 16'b0;   
     assign gt_rx_data_wire[79:64]   = 16'b0;   
     assign gt_rx_data_wire[95:80]   = 16'b0;   
     assign gt_rx_data_wire[111:96]  = 16'b0;   
     assign gt_rx_data_wire[127:112] = 16'b0; 
     assign gt_rx_data_wire[143:128] = 16'b0; 
     assign gt_rx_data_wire[159:144] = 16'b0; 
     assign gt_rx_data_wire[175:160] = 16'b0; 
     assign gt_rx_data_wire[191:176] = 16'b0; 
     assign gt_rx_data_wire[207:192] = 16'b0; 
     assign gt_rx_data_wire[223:208] = 16'b0; 
     assign gt_rx_data_wire[239:224] = 16'b0; 
     assign gt_rx_data_wire[255:240] = 16'b0; 

   end // rx_link_width_x1
  else if (LINK_CAP_MAX_LINK_WIDTH == 2)
   begin : rx_link_width_x2

     assign pipe_rx0_char_is_k =  {gt_rx_data_k_wire[1], gt_rx_data_k_wire[0]};
     assign pipe_rx1_char_is_k =  {gt_rx_data_k_wire[5], gt_rx_data_k_wire[4]};
     assign pipe_rx2_char_is_k =  2'b0 ;
     assign pipe_rx3_char_is_k =  2'b0 ;
     assign pipe_rx4_char_is_k =  2'b0 ;
     assign pipe_rx5_char_is_k =  2'b0 ;
     assign pipe_rx6_char_is_k =  2'b0 ;
     assign pipe_rx7_char_is_k =  2'b0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_k_wire[3:2]   = 2'b0; 
     assign gt_rx_data_k_wire[7:6]   = 2'b0; 
     assign gt_rx_data_k_wire[9:8]   = 2'b0; 
     assign gt_rx_data_k_wire[11:10] = 2'b0; 
     assign gt_rx_data_k_wire[13:12] = 2'b0; 
     assign gt_rx_data_k_wire[15:14] = 2'b0; 
     assign gt_rx_data_k_wire[17:16] = 2'b0; 
     assign gt_rx_data_k_wire[19:18] = 2'b0; 
     assign gt_rx_data_k_wire[21:20] = 2'b0; 
     assign gt_rx_data_k_wire[23:22] = 2'b0; 
     assign gt_rx_data_k_wire[25:24] = 2'b0; 
     assign gt_rx_data_k_wire[27:26] = 2'b0; 
     assign gt_rx_data_k_wire[29:28] = 2'b0; 
     assign gt_rx_data_k_wire[31:30] = 2'b0; 

     assign pipe_rx0_data = {gt_rx_data_wire[15: 8], gt_rx_data_wire[ 7: 0]};
     assign pipe_rx1_data = {gt_rx_data_wire[47:40], gt_rx_data_wire[39:32]} ;
     assign pipe_rx2_data = 16'h0 ;
     assign pipe_rx3_data = 16'h0 ;
     assign pipe_rx4_data = 16'h0 ;
     assign pipe_rx5_data = 16'h0 ;
     assign pipe_rx6_data = 16'h0 ;
     assign pipe_rx7_data = 16'h0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_wire[31:16]   = 16'b0; 
     assign gt_rx_data_wire[63:48]   = 16'b0;   
     assign gt_rx_data_wire[79:64]   = 16'b0;   
     assign gt_rx_data_wire[95:80]   = 16'b0;   
     assign gt_rx_data_wire[111:96]  = 16'b0;   
     assign gt_rx_data_wire[127:112] = 16'b0; 
     assign gt_rx_data_wire[143:128] = 16'b0; 
     assign gt_rx_data_wire[159:144] = 16'b0; 
     assign gt_rx_data_wire[175:160] = 16'b0; 
     assign gt_rx_data_wire[191:176] = 16'b0; 
     assign gt_rx_data_wire[207:192] = 16'b0; 
     assign gt_rx_data_wire[223:208] = 16'b0; 
     assign gt_rx_data_wire[239:224] = 16'b0; 
     assign gt_rx_data_wire[255:240] = 16'b0; 

   end // rx_link_width_x2
  else if (LINK_CAP_MAX_LINK_WIDTH == 4)
   begin : rx_link_width_x4

     assign pipe_rx0_char_is_k =  {gt_rx_data_k_wire[1], gt_rx_data_k_wire[0]};
     assign pipe_rx1_char_is_k =  {gt_rx_data_k_wire[5], gt_rx_data_k_wire[4]};
     assign pipe_rx2_char_is_k =  {gt_rx_data_k_wire[9], gt_rx_data_k_wire[8]};
     assign pipe_rx3_char_is_k =  {gt_rx_data_k_wire[13], gt_rx_data_k_wire[12]};
     assign pipe_rx4_char_is_k =  2'b0 ;
     assign pipe_rx5_char_is_k =  2'b0 ;
     assign pipe_rx6_char_is_k =  2'b0 ;
     assign pipe_rx7_char_is_k =  2'b0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_k_wire[3:2]   = 2'b0; 
     assign gt_rx_data_k_wire[7:6]   = 2'b0; 
     assign gt_rx_data_k_wire[11:10] = 2'b0; 
     assign gt_rx_data_k_wire[15:14] = 2'b0; 
     assign gt_rx_data_k_wire[17:16] = 2'b0; 
     assign gt_rx_data_k_wire[19:18] = 2'b0; 
     assign gt_rx_data_k_wire[21:20] = 2'b0; 
     assign gt_rx_data_k_wire[23:22] = 2'b0; 
     assign gt_rx_data_k_wire[25:24] = 2'b0; 
     assign gt_rx_data_k_wire[27:26] = 2'b0; 
     assign gt_rx_data_k_wire[29:28] = 2'b0; 
     assign gt_rx_data_k_wire[31:30] = 2'b0; 

     assign pipe_rx0_data = {gt_rx_data_wire[15: 8], gt_rx_data_wire[ 7: 0]};
     assign pipe_rx1_data = {gt_rx_data_wire[47:40], gt_rx_data_wire[39:32]};
     assign pipe_rx2_data = {gt_rx_data_wire[79:72], gt_rx_data_wire[71:64]};
     assign pipe_rx3_data = {gt_rx_data_wire[111:104], gt_rx_data_wire[103:96]};
     assign pipe_rx4_data = 16'h0 ;
     assign pipe_rx5_data = 16'h0 ;
     assign pipe_rx6_data = 16'h0 ;
     assign pipe_rx7_data = 16'h0 ;

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_wire[31:16]   = 16'b0; 
     assign gt_rx_data_wire[63:48]   = 16'b0;   
     assign gt_rx_data_wire[95:80]   = 16'b0;   
     assign gt_rx_data_wire[127:112] = 16'b0; 
     assign gt_rx_data_wire[143:128] = 16'b0; 
     assign gt_rx_data_wire[159:144] = 16'b0; 
     assign gt_rx_data_wire[175:160] = 16'b0; 
     assign gt_rx_data_wire[191:176] = 16'b0; 
     assign gt_rx_data_wire[207:192] = 16'b0; 
     assign gt_rx_data_wire[223:208] = 16'b0; 
     assign gt_rx_data_wire[239:224] = 16'b0; 
     assign gt_rx_data_wire[255:240] = 16'b0; 

  end // rx_link_width_x4
  else 
   begin : rx_link_width_x8

     assign pipe_rx0_char_is_k =  {gt_rx_data_k_wire[1], gt_rx_data_k_wire[0]};
     assign pipe_rx1_char_is_k =  {gt_rx_data_k_wire[5], gt_rx_data_k_wire[4]};
     assign pipe_rx2_char_is_k =  {gt_rx_data_k_wire[9], gt_rx_data_k_wire[8]};
     assign pipe_rx3_char_is_k =  {gt_rx_data_k_wire[13], gt_rx_data_k_wire[12]};
     assign pipe_rx4_char_is_k =  {gt_rx_data_k_wire[17], gt_rx_data_k_wire[16]};
     assign pipe_rx5_char_is_k =  {gt_rx_data_k_wire[21], gt_rx_data_k_wire[20]};
     assign pipe_rx6_char_is_k =  {gt_rx_data_k_wire[25], gt_rx_data_k_wire[24]};
     assign pipe_rx7_char_is_k =  {gt_rx_data_k_wire[29], gt_rx_data_k_wire[28]};

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_k_wire[3:2]   = 2'b0; 
     assign gt_rx_data_k_wire[7:6]   = 2'b0; 
     assign gt_rx_data_k_wire[11:10] = 2'b0; 
     assign gt_rx_data_k_wire[15:14] = 2'b0; 
     assign gt_rx_data_k_wire[19:18] = 2'b0; 
     assign gt_rx_data_k_wire[23:22] = 2'b0; 
     assign gt_rx_data_k_wire[27:26] = 2'b0; 
     assign gt_rx_data_k_wire[31:30] = 2'b0; 

     assign pipe_rx0_data = {gt_rx_data_wire[15: 8], gt_rx_data_wire[ 7: 0]};
     assign pipe_rx1_data = {gt_rx_data_wire[47:40], gt_rx_data_wire[39:32]};
     assign pipe_rx2_data = {gt_rx_data_wire[79:72], gt_rx_data_wire[71:64]};
     assign pipe_rx3_data = {gt_rx_data_wire[111:104], gt_rx_data_wire[103:96]};
     assign pipe_rx4_data = {gt_rx_data_wire[143:136], gt_rx_data_wire[135:128]};
     assign pipe_rx5_data = {gt_rx_data_wire[175:168], gt_rx_data_wire[167:160]};
     assign pipe_rx6_data = {gt_rx_data_wire[207:200], gt_rx_data_wire[199:192]};
     assign pipe_rx7_data = {gt_rx_data_wire[239:232], gt_rx_data_wire[231:224]};

     //synthesis warning solved: for nets below does not have driver; --assigned remaining bits of net gt_rx_data_wire to '0'
     assign gt_rx_data_wire[31:16]   = 16'b0; 
     assign gt_rx_data_wire[63:48]   = 16'b0;   
     assign gt_rx_data_wire[95:80]   = 16'b0;   
     assign gt_rx_data_wire[127:112] = 16'b0; 
     assign gt_rx_data_wire[159:144] = 16'b0; 
     assign gt_rx_data_wire[191:176] = 16'b0; 
     assign gt_rx_data_wire[223:208] = 16'b0; 
     assign gt_rx_data_wire[255:240] = 16'b0; 

  end // rx_link_width_x8
endgenerate

assign pipe_rx0_status = gt_rx_status_wire[ 2: 0];
assign pipe_rx1_status = (LINK_CAP_MAX_LINK_WIDTH >= 2 ) ? gt_rx_status_wire[ 5: 3] : 3'b0 ;
assign pipe_rx2_status = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_status_wire[ 8: 6] : 3'b0 ;
assign pipe_rx3_status = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_status_wire[11: 9] : 3'b0 ;
assign pipe_rx4_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_status_wire[14:12] : 3'b0 ;
assign pipe_rx5_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_status_wire[17:15] : 3'b0 ;
assign pipe_rx6_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_status_wire[20:18] : 3'b0 ;
assign pipe_rx7_status = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_status_wire[23:21] : 3'b0 ;

//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<
//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<

assign pipe_rx0_elec_idle = gt_rx_elec_idle_wire[0];
assign pipe_rx1_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 2 ) ? gt_rx_elec_idle_wire[1] : 1'b1 ;
assign pipe_rx2_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_elec_idle_wire[2] : 1'b1 ;
assign pipe_rx3_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_elec_idle_wire[3] : 1'b1 ;
assign pipe_rx4_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_elec_idle_wire[4] : 1'b1 ;
assign pipe_rx5_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_elec_idle_wire[5] : 1'b1 ;
assign pipe_rx6_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_elec_idle_wire[6] : 1'b1 ;
assign pipe_rx7_elec_idle = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_elec_idle_wire[7] : 1'b1 ;

assign pipe_rx0_valid = gt_rx_valid_wire[0];
assign pipe_rx1_valid = (LINK_CAP_MAX_LINK_WIDTH >= 2 ) ? gt_rx_valid_wire[1] : 1'b0 ;
assign pipe_rx2_valid = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_valid_wire[2] : 1'b0 ;
assign pipe_rx3_valid = (LINK_CAP_MAX_LINK_WIDTH >= 4 ) ? gt_rx_valid_wire[3] : 1'b0 ;
assign pipe_rx4_valid = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_valid_wire[4] : 1'b0 ;
assign pipe_rx5_valid = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_valid_wire[5] : 1'b0 ;
assign pipe_rx6_valid = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_valid_wire[6] : 1'b0 ;
assign pipe_rx7_valid = (LINK_CAP_MAX_LINK_WIDTH >= 8 ) ? gt_rx_valid_wire[7] : 1'b0 ;

assign gt_rx_polarity[0] = pipe_rx0_polarity;
assign gt_rx_polarity[1] = pipe_rx1_polarity;
assign gt_rx_polarity[2] = pipe_rx2_polarity;
assign gt_rx_polarity[3] = pipe_rx3_polarity;
assign gt_rx_polarity[4] = pipe_rx4_polarity;
assign gt_rx_polarity[5] = pipe_rx5_polarity;
assign gt_rx_polarity[6] = pipe_rx6_polarity;
assign gt_rx_polarity[7] = pipe_rx7_polarity;

assign gt_power_down[ 1: 0] = pipe_tx0_powerdown;
assign gt_power_down[ 3: 2] = pipe_tx1_powerdown;
assign gt_power_down[ 5: 4] = pipe_tx2_powerdown;
assign gt_power_down[ 7: 6] = pipe_tx3_powerdown;
assign gt_power_down[ 9: 8] = pipe_tx4_powerdown;
assign gt_power_down[11:10] = pipe_tx5_powerdown;
assign gt_power_down[13:12] = pipe_tx6_powerdown;
assign gt_power_down[15:14] = pipe_tx7_powerdown;

assign gt_tx_char_disp_mode = {pipe_tx7_compliance,
                               pipe_tx6_compliance,
                               pipe_tx5_compliance,
                               pipe_tx4_compliance,
                               pipe_tx3_compliance,
                               pipe_tx2_compliance,
                               pipe_tx1_compliance,
                               pipe_tx0_compliance};


assign gt_tx_data_k = {2'd0,
                       pipe_tx7_char_is_k,
                       2'd0,
                       pipe_tx6_char_is_k,
                       2'd0,
                       pipe_tx5_char_is_k,
                       2'd0,
                       pipe_tx4_char_is_k,
                       2'd0,
                       pipe_tx3_char_is_k,
                       2'd0,
                       pipe_tx2_char_is_k,
                       2'd0,
                       pipe_tx1_char_is_k,
                       2'd0,
                       pipe_tx0_char_is_k};

assign gt_tx_data = {16'd0,
                     pipe_tx7_data,
                     16'd0,
                     pipe_tx6_data,
                     16'd0,
                     pipe_tx5_data,
                     16'd0,
                     pipe_tx4_data,
                     16'd0,
                     pipe_tx3_data,
                     16'd0,
                     pipe_tx2_data,
                     16'd0,
                     pipe_tx1_data,
                     16'd0,
                     pipe_tx0_data};

assign gt_tx_detect_rx_loopback = pipe_tx_rcvr_det;

assign gt_tx_elec_idle = {pipe_tx7_elec_idle,
                          pipe_tx6_elec_idle,
                          pipe_tx5_elec_idle,
                          pipe_tx4_elec_idle,
                          pipe_tx3_elec_idle,
                          pipe_tx2_elec_idle,
                          pipe_tx1_elec_idle,
                          pipe_tx0_elec_idle};

always @(posedge pipe_clk_int or negedge clock_locked) begin
  if (!clock_locked)
    reg_clock_locked <= #TCQ 1'b0;
  else
    reg_clock_locked <= #TCQ 1'b1;
end

always @(posedge pipe_clk_int) begin
  if (!reg_clock_locked)
    phy_rdy_n_int <= #TCQ 1'b0;
  else
    phy_rdy_n_int <= #TCQ all_phystatus_rst;
end

assign all_phystatus_rst = (&phystatus_rst[LINK_CAP_MAX_LINK_WIDTH-1:0]);
assign phy_rdy_n     = phy_rdy_n_int;

endmodule


`timescale 1ns/1ps
module model_ap2_tst_gt_rx_valid_filter_7x #(

  parameter           CLK_COR_MIN_LAT    = 28,
  parameter           TCQ                = 1

)
(
  output  [1:0]       USER_RXCHARISK,
  output  [15:0]      USER_RXDATA,
  output              USER_RXVALID,
  output              USER_RXELECIDLE,
  output  [ 2:0]      USER_RX_STATUS,
  output              USER_RX_PHY_STATUS,
  input  [1:0]        GT_RXCHARISK,
  input  [15:0]       GT_RXDATA,
  input               GT_RXVALID,
  input               GT_RXELECIDLE,
  input  [ 2:0]       GT_RX_STATUS,
  input               GT_RX_PHY_STATUS,

  input               PLM_IN_L0,
  input               PLM_IN_RS,

  input               USER_CLK,
  input               RESET

);



  localparam EIOS_DET_IDL      = 5'b00001;
  localparam EIOS_DET_NO_STR0  = 5'b00010;
  localparam EIOS_DET_STR0     = 5'b00100;
  localparam EIOS_DET_STR1     = 5'b01000;
  localparam EIOS_DET_DONE     = 5'b10000;

  localparam EIOS_COM          = 8'hBC;
  localparam EIOS_IDL          = 8'h7C;
  localparam FTSOS_COM         = 8'hBC;
  localparam FTSOS_FTS         = 8'h3C;

  reg    [4:0]        reg_state_eios_det;
  wire   [4:0]        state_eios_det;

  reg                 reg_eios_detected;
  wire                eios_detected;

  reg                 reg_symbol_after_eios;
  wire                symbol_after_eios;

  localparam USER_RXVLD_IDL     = 4'b0001;
  localparam USER_RXVLD_EI      = 4'b0010;
  localparam USER_RXVLD_EI_DB0  = 4'b0100;
  localparam USER_RXVLD_EI_DB1  = 4'b1000;


  reg    [1:0]        gt_rxcharisk_q;
  reg    [15:0]       gt_rxdata_q;
  reg                 gt_rxvalid_q;
  reg                 gt_rxelecidle_q;

  reg    [ 2:0]       gt_rx_status_q;
  reg                 gt_rx_phy_status_q;
  reg                 gt_rx_is_skp0_q;
  reg                 gt_rx_is_skp1_q;

  // EIOS detector

  always @(posedge USER_CLK) begin

    if (RESET) begin

      reg_eios_detected <= #TCQ 1'b0;
      reg_state_eios_det <= #TCQ EIOS_DET_IDL;
      reg_symbol_after_eios <= #TCQ 1'b0;
      gt_rxcharisk_q <= #TCQ 2'b00;
      gt_rxdata_q <= #TCQ 16'h0;
      gt_rxvalid_q <= #TCQ 1'b0;
      gt_rxelecidle_q <= #TCQ 1'b0;
      gt_rx_status_q <= #TCQ 3'b000;
      gt_rx_phy_status_q <= #TCQ 1'b0;
      gt_rx_is_skp0_q <= #TCQ 1'b0;
      gt_rx_is_skp1_q <= #TCQ 1'b0;

    end else begin
      reg_eios_detected <= #TCQ 1'b0;
      reg_symbol_after_eios <= #TCQ 1'b0;
        gt_rxcharisk_q <= #TCQ GT_RXCHARISK;
        gt_rxelecidle_q <= #TCQ GT_RXELECIDLE;
      gt_rxdata_q <= #TCQ GT_RXDATA;
      gt_rx_phy_status_q <= #TCQ GT_RX_PHY_STATUS;
      
     //De-assert rx_valid signal when EIOS is detected on RXDATA
      if(((reg_state_eios_det == 5'b10000)) && (PLM_IN_L0)
       ) begin
       
        gt_rxvalid_q <= #TCQ 1'b0; 
      end
      else if (GT_RXELECIDLE && !gt_rxvalid_q) begin
         gt_rxvalid_q <= #TCQ 1'b0; 
      end   
      else begin
       gt_rxvalid_q <= GT_RXVALID;
     end  

     if (gt_rxvalid_q) begin
      gt_rx_status_q <= #TCQ GT_RX_STATUS;
       
     end
     else if (!gt_rxvalid_q && PLM_IN_L0) begin
      gt_rx_status_q <= #TCQ 3'b0;
     end
     else begin
      gt_rx_status_q <= #TCQ GT_RX_STATUS;
     end  

      
      
      if (GT_RXCHARISK[0] && GT_RXDATA[7:0] == FTSOS_FTS)
        gt_rx_is_skp0_q <= #TCQ 1'b1;
      else
        gt_rx_is_skp0_q <= #TCQ 1'b0;

      if (GT_RXCHARISK[1] && GT_RXDATA[15:8] == FTSOS_FTS)
        gt_rx_is_skp1_q <= #TCQ 1'b1;
      else
        gt_rx_is_skp1_q <= #TCQ 1'b0;

      case ( state_eios_det )

        EIOS_DET_IDL : begin

          if ((gt_rxcharisk_q[0]) && (gt_rxdata_q[7:0] == EIOS_COM) &&
              (gt_rxcharisk_q[1]) && (gt_rxdata_q[15:8] == EIOS_IDL)) begin

            reg_state_eios_det <= #TCQ EIOS_DET_NO_STR0;
            reg_eios_detected <= #TCQ 1'b1;
          //  gt_rxvalid_q <= #TCQ 1'b0;

          end else if ((gt_rxcharisk_q[1]) && (gt_rxdata_q[15:8] == EIOS_COM))
            reg_state_eios_det <= #TCQ EIOS_DET_STR0;
          else
            reg_state_eios_det <= #TCQ EIOS_DET_IDL;

        end

        EIOS_DET_NO_STR0 : begin

          if ((gt_rxcharisk_q[0] && (gt_rxdata_q[7:0] == EIOS_IDL)) &&
              (gt_rxcharisk_q[1] && (gt_rxdata_q[15:8] == EIOS_IDL)))
              begin
            reg_state_eios_det <= #TCQ EIOS_DET_DONE;
            gt_rxvalid_q <= #TCQ 1'b0;
            end
         else if (gt_rxcharisk_q[0] && (gt_rxdata_q[7:0] == EIOS_IDL)) begin
            
            reg_state_eios_det <= #TCQ EIOS_DET_DONE;
            gt_rxvalid_q <= #TCQ 1'b0;
            end
          else
            reg_state_eios_det <= #TCQ EIOS_DET_IDL;

        end

        EIOS_DET_STR0 : begin

          if ((gt_rxcharisk_q[0] && (gt_rxdata_q[7:0] == EIOS_IDL)) &&
              (gt_rxcharisk_q[1] && (gt_rxdata_q[15:8] == EIOS_IDL))) begin

            reg_state_eios_det <= #TCQ EIOS_DET_STR1;
            reg_eios_detected <= #TCQ 1'b1;
            gt_rxvalid_q <= #TCQ 1'b0;
            reg_symbol_after_eios <= #TCQ 1'b1;

          end else
            reg_state_eios_det <= #TCQ EIOS_DET_IDL;

        end

        EIOS_DET_STR1 : begin

          if ((gt_rxcharisk_q[0]) && (gt_rxdata_q[7:0] == EIOS_IDL))
          begin
            reg_state_eios_det <= #TCQ EIOS_DET_DONE;
            gt_rxvalid_q <= #TCQ 1'b0;
          end  
          else
            reg_state_eios_det <= #TCQ EIOS_DET_IDL;

        end

        EIOS_DET_DONE : begin

          reg_state_eios_det <= #TCQ EIOS_DET_IDL;

        end

      endcase

    end

  end
  assign state_eios_det = reg_state_eios_det;
  assign eios_detected = reg_eios_detected;
  assign symbol_after_eios = reg_symbol_after_eios;
  /*SRL16E #(.INIT(0)) rx_elec_idle_delay (.Q(USER_RXELECIDLE),
                                         .D(gt_rxelecidle_q),
                                         .CLK(USER_CLK),
                                         .CE(1'b1), .A3(1'b1),.A2(1'b1),.A1(1'b1),.A0(1'b1));
*/
wire    rst_l = ~RESET;


assign USER_RXVALID = gt_rxvalid_q;
assign USER_RXCHARISK[0] = gt_rxvalid_q ? gt_rxcharisk_q[0] : 1'b0;
assign USER_RXCHARISK[1] = (gt_rxvalid_q && !symbol_after_eios) ? gt_rxcharisk_q[1] : 1'b0;
assign USER_RXDATA[7:0] = gt_rxdata_q[7:0];
assign USER_RXDATA[15:8] = gt_rxdata_q[15:8];
assign USER_RX_STATUS = gt_rx_status_q;
assign USER_RX_PHY_STATUS = gt_rx_phy_status_q;
assign USER_RXELECIDLE = gt_rxelecidle_q;


endmodule


`timescale 1ns/1ps
module model_ap2_tst_pipe_wrapper #
(

    parameter PCIE_SIM_MODE                 = "FALSE",      // PCIe sim mode 
    parameter PCIE_SIM_SPEEDUP              = "FALSE",      // PCIe sim speedup
    parameter PCIE_SIM_TX_EIDLE_DRIVE_LEVEL = "1",          // PCIe sim TX electrical idle drive level 
    parameter PCIE_GT_DEVICE                = "GTX",        // PCIe GT device
    parameter PCIE_USE_MODE                 = "3.0",        // PCIe use mode
    parameter PCIE_PLL_SEL                  = "CPLL",       // PCIe PLL select for Gen1/Gen2 (GTX/GTH) only
    parameter PCIE_AUX_CDR_GEN3_EN          = "TRUE",       // PCIe AUX CDR for Gen3 (GTH 2.0) only
    parameter PCIE_LPM_DFE                  = "LPM",        // PCIe LPM or DFE mode for Gen1/Gen2 only
    parameter PCIE_LPM_DFE_GEN3             = "DFE",        // PCIe LPM or DFE mode for Gen3      only
    parameter PCIE_EXT_CLK                  = "FALSE",      // PCIe external clock
    parameter PCIE_EXT_GT_COMMON            = "FALSE",      // PCIe external GT COMMON
    parameter EXT_CH_GT_DRP                 = "FALSE",      // PCIe external CH DRP

    parameter TX_MARGIN_FULL_0              = 7'b1001111,                          // 1000 mV
    parameter TX_MARGIN_FULL_1              = 7'b1001110,                          // 950 mV
    parameter TX_MARGIN_FULL_2              = 7'b1001101,                          // 900 mV
    parameter TX_MARGIN_FULL_3              = 7'b1001100,                          // 850 mV
    parameter TX_MARGIN_FULL_4              = 7'b1000011,                          // 400 mV
    parameter TX_MARGIN_LOW_0               = 7'b1000101,                          // 500 mV
    parameter TX_MARGIN_LOW_1               = 7'b1000110 ,                          // 450 mV
    parameter TX_MARGIN_LOW_2               = 7'b1000011,                          // 400 mV
    parameter TX_MARGIN_LOW_3               = 7'b1000010 ,                          // 350 mV
    parameter TX_MARGIN_LOW_4               = 7'b1000000 ,

    parameter PCIE_POWER_SAVING             = "TRUE",       // PCIe power saving
    parameter PCIE_ASYNC_EN                 = "FALSE",      // PCIe async enable
    parameter PCIE_TXBUF_EN                 = "FALSE",      // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_RXBUF_EN                 = "TRUE",       // PCIe RX buffer enable for Gen3      only
    parameter PCIE_TXSYNC_MODE              = 0,            // PCIe TX sync mode
    parameter PCIE_RXSYNC_MODE              = 0,            // PCIe RX sync mode
    parameter PCIE_CHAN_BOND                = 1,            // PCIe channel bonding mode
    parameter PCIE_CHAN_BOND_EN             = "TRUE",       // PCIe channel bonding enable for Gen1/Gen2 only
    parameter PCIE_LANE                     = 1,            // PCIe number of lanes
    parameter PCIE_LINK_SPEED               = 3,            // PCIe link speed 
    parameter PCIE_REFCLK_FREQ              = 0,            // PCIe reference clock frequency
    parameter PCIE_USERCLK1_FREQ            = 2,            // PCIe user clock 1 frequency
    parameter PCIE_USERCLK2_FREQ            = 2,            // PCIe user clock 2 frequency
    parameter PCIE_TX_EIDLE_ASSERT_DELAY    = 3'd4,         // PCIe TX electrical idle assert delay
    parameter PCIE_RXEQ_MODE_GEN3           = 1,            // PCIe RX equalization mode
    parameter PCIE_OOBCLK_MODE              = 1,            // PCIe OOB clock mode
    parameter PCIE_JTAG_MODE                = 0,            // PCIe JTAG mode
    parameter PCIE_DEBUG_MODE               = 0             // PCIe debug mode 
    
)                                                     
                                                            //--------------------------------------
(                                                           // Gen1/Gen2  | Gen3 
                                                            //--------------------------------------
    //---------- PIPE Clock & Reset Ports ------------------
    input                           PIPE_CLK,               // Reference clock that drives MMCM
    input                           PIPE_RESET_N,           // PCLK       | PCLK
   
    output                          PIPE_PCLK,              // Drives [TX/RX]USRCLK in Gen1/Gen2
                                                            // Drives TXUSRCLK in Gen3
                                                            // Drives RXUSRCLK in Gen3 async mode only
    //---------- PIPE TX Data Ports ------------------------
    input       [(PCIE_LANE*32)-1:0]PIPE_TXDATA,            // PCLK       | PCLK
    input       [(PCIE_LANE*4)-1:0] PIPE_TXDATAK,           // PCLK       | PCLK
    
    output      [PCIE_LANE-1:0]     PIPE_TXP,               // Serial data
    output      [PCIE_LANE-1:0]     PIPE_TXN,               // Serial data

    //---------- PIPE RX Data Ports ------------------------
    input       [PCIE_LANE-1:0]     PIPE_RXP,               // Serial data
    input       [PCIE_LANE-1:0]     PIPE_RXN,               // Serial data
    
    output      [(PCIE_LANE*32)-1:0]PIPE_RXDATA,            // PCLK       | RXUSRCLK
    output      [(PCIE_LANE*4)-1:0] PIPE_RXDATAK,           // PCLK       | RXUSRCLK
    
    //---------- PIPE Command Ports ------------------------
    input                           PIPE_TXDETECTRX,        // PCLK       | PCLK
    input       [PCIE_LANE-1:0]     PIPE_TXELECIDLE,        // PCLK       | PCLK
    input       [PCIE_LANE-1:0]     PIPE_TXCOMPLIANCE,      // PCLK       | PCLK   
    input       [PCIE_LANE-1:0]     PIPE_RXPOLARITY,        // PCLK       | RXUSRCLK
    input       [(PCIE_LANE*2)-1:0] PIPE_POWERDOWN,         // PCLK       | PCLK
    input       [ 1:0]              PIPE_RATE,              // PCLK       | PCLK
    
    //---------- PIPE Electrical Command Ports -------------   
    input       [ 2:0]              PIPE_TXMARGIN,          // Async      | Async 
    input                           PIPE_TXSWING,           // Async      | Async 
    input       [PCIE_LANE-1:0]     PIPE_TXDEEMPH,          // Async/PCLK | Async/PCLK  
    input       [(PCIE_LANE*2)-1:0] PIPE_TXEQ_CONTROL,      // PCLK       | PCLK  
    input       [(PCIE_LANE*4)-1:0] PIPE_TXEQ_PRESET,       // PCLK       | PCLK  
    input       [(PCIE_LANE*4)-1:0] PIPE_TXEQ_PRESET_DEFAULT,// PCLK      | PCLK 
    input       [(PCIE_LANE*6)-1:0] PIPE_TXEQ_DEEMPH,       // PCLK       | PCLK  
                                                                            
    input       [(PCIE_LANE*2)-1:0] PIPE_RXEQ_CONTROL,      // PCLK       | PCLK  
    input       [(PCIE_LANE*3)-1:0] PIPE_RXEQ_PRESET,       // PCLK       | PCLK  
    input       [(PCIE_LANE*6)-1:0] PIPE_RXEQ_LFFS,         // PCLK       | PCLK  
    input       [(PCIE_LANE*4)-1:0] PIPE_RXEQ_TXPRESET,     // PCLK       | PCLK  
    input       [PCIE_LANE-1:0]     PIPE_RXEQ_USER_EN,      // PCLK       | PCLK      
    input       [(PCIE_LANE*18)-1:0]PIPE_RXEQ_USER_TXCOEFF, // PCLK       | PCLK
    input       [PCIE_LANE-1:0]     PIPE_RXEQ_USER_MODE,    // PCLK       | PCLK
                                                                           
    output      [ 5:0]              PIPE_TXEQ_FS,           // Async      | Async  
    output      [ 5:0]              PIPE_TXEQ_LF,           // Async      | Async 
    output      [(PCIE_LANE*18)-1:0]PIPE_TXEQ_COEFF,        // PCLK       | PCLK  
    output      [PCIE_LANE-1:0]     PIPE_TXEQ_DONE,         // PCLK       | PCLK  
                                                                           
    output      [(PCIE_LANE*18)-1:0]PIPE_RXEQ_NEW_TXCOEFF,  // PCLK       | PCLK  
    output      [PCIE_LANE-1:0]     PIPE_RXEQ_LFFS_SEL,     // PCLK       | PCLK  
    output      [PCIE_LANE-1:0]     PIPE_RXEQ_ADAPT_DONE,   // PCLK       | PCLK  
    output      [PCIE_LANE-1:0]     PIPE_RXEQ_DONE,         // PCLK       | PCLK  
    
    //---------- PIPE Status Ports -------------------------
    output      [PCIE_LANE-1:0]     PIPE_RXVALID,           // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_PHYSTATUS,         // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_PHYSTATUS_RST,     // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_RXELECIDLE,        // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_EYESCANDATAERROR,  // Async      | Async
    output      [(PCIE_LANE*3)-1:0] PIPE_RXSTATUS,          // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_RXPMARESETDONE,    // Async      | Async
    output      [(PCIE_LANE*3)-1:0] PIPE_RXBUFSTATUS,       // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_TXPHALIGNDONE,     // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_TXPHINITDONE,      // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_TXDLYSRESETDONE,   // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_RXPHALIGNDONE,     // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_RXDLYSRESETDONE,   // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_RXSYNCDONE,        // PCLK       | RXUSRCLK
    output      [(PCIE_LANE*8)-1:0] PIPE_RXDISPERR,         // PCLK       | RXUSRCLK
    output      [(PCIE_LANE*8)-1:0] PIPE_RXNOTINTABLE,      // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_RXCOMMADET,        // PCLK       | RXUSRCLK
    
    //---------- PIPE User Ports ---------------------------
    input                           PIPE_MMCM_RST_N,        // Async      | Async
    input       [PCIE_LANE-1:0]     PIPE_RXSLIDE,           // PCLK       | RXUSRCLK
    
    output      [PCIE_LANE-1:0]     PIPE_CPLL_LOCK,         // Async      | Async
    output      [(PCIE_LANE-1)>>2:0]PIPE_QPLL_LOCK,         // Async      | Async
    output                          PIPE_PCLK_LOCK,         // Async      | Async
    output      [PCIE_LANE-1:0]     PIPE_RXCDRLOCK,         // Async      | Async
    output                          PIPE_USERCLK1,          // Optional user clock
    output                          PIPE_USERCLK2,          // Optional user clock
    output                          PIPE_RXUSRCLK,          // RXUSRCLK 
                                                            // Equivalent to PCLK in Gen1/Gen2
                                                            // Equivalent to RXOUTCLK[0] in Gen3
    output      [PCIE_LANE-1:0]     PIPE_RXOUTCLK,          // RX recovered clock (for debug only)
    output      [PCIE_LANE-1:0]     PIPE_TXSYNC_DONE,       // PCLK       | PCLK
    output      [PCIE_LANE-1:0]     PIPE_RXSYNC_DONE,       // PCLK       | PCLK
    output      [PCIE_LANE-1:0]     PIPE_GEN3_RDY,          // PCLK       | RXUSRCLK
    output      [PCIE_LANE-1:0]     PIPE_RXCHANISALIGNED,
    output      [PCIE_LANE-1:0]     PIPE_ACTIVE_LANE,

// Shared Logic Internal
    output                          INT_PCLK_OUT_SLAVE,     // PCLK       | PCLK
    output                          INT_RXUSRCLK_OUT,       // RXUSERCLK
    output  [PCIE_LANE-1:0  ]       INT_RXOUTCLK_OUT,       // RX recovered clock
    output                          INT_DCLK_OUT,           // DCLK       | DCLK
    output                          INT_USERCLK1_OUT,       // Optional user clock
    output                          INT_USERCLK2_OUT,       // Optional user clock
    output                          INT_OOBCLK_OUT,         // OOB        | OOB
    output                          INT_MMCM_LOCK_OUT,      // Async      | Async
    output  [1:0]                   INT_QPLLLOCK_OUT,
    output  [1:0]                   INT_QPLLOUTCLK_OUT,
    output  [1:0]                   INT_QPLLOUTREFCLK_OUT,
    input   [PCIE_LANE-1:0]         INT_PCLK_SEL_SLAVE,

  // Shared Logic External
    
    //---------- External Clock Ports ----------------------
    input                           PIPE_PCLK_IN,           // PCLK       | PCLK
    input                           PIPE_RXUSRCLK_IN,       // RXUSERCLK
                                                            // Equivalent to PCLK in Gen1/Gen2
                                                            // Equivalent to RXOUTCLK[0] in Gen3
    input       [PCIE_LANE-1:0]     PIPE_RXOUTCLK_IN,       // RX recovered clock
    input                           PIPE_DCLK_IN,           // DCLK       | DCLK
    input                           PIPE_USERCLK1_IN,       // Optional user clock
    input                           PIPE_USERCLK2_IN,       // Optional user clock
    input                           PIPE_OOBCLK_IN,         // OOB        | OOB
    input                           PIPE_MMCM_LOCK_IN,      // Async      | Async
    
    output                          PIPE_TXOUTCLK_OUT,      // PCLK       | PCLK
    output      [PCIE_LANE-1:0]     PIPE_RXOUTCLK_OUT,      // RX recovered clock (for debug only)
    output      [PCIE_LANE-1:0]     PIPE_PCLK_SEL_OUT,      // PCLK       | PCLK
    output                          PIPE_GEN3_OUT,          // PCLK       | PCLK
    //---------- External GT COMMON Ports ----------------------
    input       [11:0]              QPLL_DRP_CRSCODE,
    input       [17:0]              QPLL_DRP_FSM,
    input       [1:0]               QPLL_DRP_DONE,
    input       [1:0]               QPLL_DRP_RESET,
    input       [1:0]               QPLL_QPLLLOCK,
    input       [1:0]               QPLL_QPLLOUTCLK,
    input       [1:0]               QPLL_QPLLOUTREFCLK,
    output              	          QPLL_QPLLPD,
    output      [1:0]               QPLL_QPLLRESET,
    output              	          QPLL_DRP_CLK,
    output              	          QPLL_DRP_RST_N,
    output              	          QPLL_DRP_OVRD,
    output              	          QPLL_DRP_GEN3,
    output              	          QPLL_DRP_START,

    //---------- TRANSCEIVER DEBUG -----------------------
    input       [ 2:0]              PIPE_TXPRBSSEL,         // PCLK       | PCLK
    input       [ 2:0]              PIPE_RXPRBSSEL,         // PCLK       | PCLK
    input                           PIPE_TXPRBSFORCEERR,    // PCLK       | PCLK
    input                           PIPE_RXPRBSCNTRESET,    // PCLK       | PCLK
    input       [ 2:0]              PIPE_LOOPBACK,          // PCLK       | PCLK
    
    output      [PCIE_LANE-1:0]     PIPE_RXPRBSERR,         // PCLK       | PCLK
    
    //---------- FSM Ports ---------------------------------
    output      [4:0]               PIPE_RST_FSM,           // PCLK       | PCLK
    output      [11:0]              PIPE_QRST_FSM,          // PCLK       | PCLK
    output      [(PCIE_LANE*5)-1:0] PIPE_RATE_FSM,          // PCLK       | PCLK
    output      [(PCIE_LANE*6)-1:0] PIPE_SYNC_FSM_TX,       // PCLK       | PCLK
    output      [(PCIE_LANE*7)-1:0] PIPE_SYNC_FSM_RX,       // PCLK       | PCLK
    output      [(PCIE_LANE*7)-1:0] PIPE_DRP_FSM,           // DCLK       | DCLK
    output      [(PCIE_LANE*6)-1:0] PIPE_TXEQ_FSM,          // PCLK       | PCLK
    output      [(PCIE_LANE*6)-1:0] PIPE_RXEQ_FSM,          // PCLK       | PCLK
    output      [((((PCIE_LANE-1)>>2)+1)*9)-1:0]PIPE_QDRP_FSM, // DCLK    | DCLK  
        
    output                          PIPE_RST_IDLE,          // PCLK       | PCLK 
    output                          PIPE_QRST_IDLE,         // PCLK       | PCLK 
    output                          PIPE_RATE_IDLE,         // PCLK       | PCLK 
    
    //----------- Channel DRP----------------------------
    output                            EXT_CH_GT_DRPCLK,
    input        [(PCIE_LANE*9)-1:0] EXT_CH_GT_DRPADDR,
    input        [PCIE_LANE-1:0]     EXT_CH_GT_DRPEN,
    input        [(PCIE_LANE*16)-1:0]EXT_CH_GT_DRPDI,
    input        [PCIE_LANE-1:0]     EXT_CH_GT_DRPWE,

    output       [(PCIE_LANE*16)-1:0]EXT_CH_GT_DRPDO,
    output       [PCIE_LANE-1:0]     EXT_CH_GT_DRPRDY,

    //---------- JTAG Ports --------------------------------
    input                           PIPE_JTAG_EN,           // DCLK       | DCLK
    output      [PCIE_LANE-1:0]     PIPE_JTAG_RDY,          // DCLK       | DCLK
    
    //---------- Debug Ports -------------------------------
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_0,           // Async      | Async 
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_1,           // Async      | Async 
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_2,           // Async      | Async 
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_3,           // Async      | Async 
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_4,           // Async      | Async 
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_5,           // Async      | Async   
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_6,           // Async      | Async   
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_7,           // Async      | Async   
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_8,           // Async      | Async   
    output      [PCIE_LANE-1:0]     PIPE_DEBUG_9,           // Async      | Async   
    output      [31:0]              PIPE_DEBUG,             // Async      | Async 
    
    output      [(PCIE_LANE*15)-1:0] PIPE_DMONITOROUT       // DMONITORCLK
    
);

    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             reset_n_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             reset_n_reg2;

    //---------- PIPE Clock Module Output ------------------ 
    wire                            clk_pclk;  
    wire                            clk_rxusrclk;
    wire        [PCIE_LANE-1:0]     clk_rxoutclk;
    wire                            clk_dclk;
    wire                            clk_oobclk;
    wire                            clk_mmcm_lock;
    
    //---------- PIPE Reset Module Output ------------------
    wire                            rst_cpllreset;
    wire                            rst_cpllpd;
    wire                            rst_rxusrclk_reset;
    wire                            rst_dclk_reset;   
    wire rst_gtreset;
    wire                            rst_drp_start;
    wire                            rst_drp_x16x20_mode;
    wire                            rst_drp_x16;
    wire rst_userrdy;
    wire                            rst_txsync_start;
    wire                            rst_idle;
    wire        [4:0]               rst_fsm;
    
    //------------------------------------------------------
    wire                            gtp_rst_qpllreset;      // GTP
    wire                            gtp_rst_qpllpd;         // GTP
    
    //------------------------------------------------------
    wire        [(PCIE_LANE-1)>>2:0]qpllreset;          
    wire                            qpllpd;
    
    //---------- QPLL Reset Module Output ------------------
    wire                            qrst_ovrd;
    wire                            qrst_drp_start;
    wire                            qrst_qpllreset;
    wire                            qrst_qpllpd;
    wire                            qrst_idle;
    wire        [3:0]               qrst_fsm;
    
    //---------- PIPE_JTAG Master Module Output ------------
    wire        [(PCIE_LANE*37)-1:0] jtag_sl_iport;
    wire        [(PCIE_LANE*17)-1:0] jtag_sl_oport;
    
    //---------- PIPE User Module Output -------------------
    wire [PCIE_LANE-1:0] gt_txpmareset_i;                 
    wire [PCIE_LANE-1:0] gt_rxpmareset_i;                 

    wire        [PCIE_LANE-1:0]     user_oobclk;
    wire        [PCIE_LANE-1:0]     user_resetovrd;
    wire        [PCIE_LANE-1:0]     user_txpmareset;                 
    wire        [PCIE_LANE-1:0]     user_rxpmareset;                
    wire        [PCIE_LANE-1:0]     user_rxcdrreset;
    wire        [PCIE_LANE-1:0]     user_rxcdrfreqreset;
    wire [PCIE_LANE-1:0] user_rxdfelpmreset;
    wire [PCIE_LANE-1:0] user_eyescanreset;
    wire [PCIE_LANE-1:0] user_txpcsreset;                   
    wire [PCIE_LANE-1:0] user_rxpcsreset;                 
    wire [PCIE_LANE-1:0] user_rxbufreset;
    wire        [PCIE_LANE-1:0]     user_resetovrd_done;
    wire        [PCIE_LANE-1:0]     user_active_lane;
    wire        [PCIE_LANE-1:0]     user_resetdone /* synthesis syn_keep=1 */;
    wire        [PCIE_LANE-1:0]     user_rxcdrlock;
    wire        [PCIE_LANE-1:0]     user_rx_converge; 
    wire        [PCIE_LANE-1:0]     PIPE_RXEQ_CONVERGE;
    
    //---------- PIPE Rate Module Output -------------------
    wire        [PCIE_LANE-1:0]     rate_cpllpd;
    wire        [PCIE_LANE-1:0]     rate_qpllpd;
    wire        [PCIE_LANE-1:0]     rate_cpllreset;
    wire        [PCIE_LANE-1:0]     rate_qpllreset;
    wire        [PCIE_LANE-1:0]     rate_txpmareset;
    wire        [PCIE_LANE-1:0]     rate_rxpmareset;
    wire        [(PCIE_LANE*2)-1:0] rate_sysclksel;
    wire        [PCIE_LANE-1:0]     rate_pclk_sel;
    wire        [PCIE_LANE-1:0]     rate_drp_start;
    wire        [PCIE_LANE-1:0]     rate_drp_x16x20_mode;
    wire        [PCIE_LANE-1:0]     rate_drp_x16;
    wire        [PCIE_LANE-1:0]     rate_gen3;
    wire        [(PCIE_LANE*3)-1:0] rate_rate;
    wire        [PCIE_LANE-1:0]     rate_resetovrd_start;
    wire        [PCIE_LANE-1:0]     rate_txsync_start;
    wire        [PCIE_LANE-1:0]     rate_done;
    wire        [PCIE_LANE-1:0]     rate_rxsync_start;
    wire        [PCIE_LANE-1:0]     rate_rxsync;
    wire        [PCIE_LANE-1:0]     rate_idle;
    wire        [(PCIE_LANE*5)-1:0] rate_fsm;

    //---------- PIPE Sync Module Output -------------------
    wire        [PCIE_LANE-1:0]     sync_txphdlyreset;
    wire        [PCIE_LANE-1:0]     sync_txphalign;    
    wire        [PCIE_LANE-1:0]     sync_txphalignen; 
    wire        [PCIE_LANE-1:0]     sync_txphinit;   
    wire        [PCIE_LANE-1:0]     sync_txdlybypass; 
    wire        [PCIE_LANE-1:0]     sync_txdlysreset;   
    wire        [PCIE_LANE-1:0]     sync_txdlyen;      
    wire        [PCIE_LANE-1:0]     sync_txsync_done;
    wire        [(PCIE_LANE*6)-1:0] sync_fsm_tx;
    
    wire        [PCIE_LANE-1:0]     sync_rxphalign;
    wire        [PCIE_LANE-1:0]     sync_rxphalignen;
    wire        [PCIE_LANE-1:0]     sync_rxdlybypass;
    wire        [PCIE_LANE-1:0]     sync_rxdlysreset;
    wire        [PCIE_LANE-1:0]     sync_rxdlyen;
    wire        [PCIE_LANE-1:0]     sync_rxddien;
    wire        [PCIE_LANE-1:0]     sync_rxsync_done; 
    wire        [PCIE_LANE-1:0]     sync_rxsync_donem;      
    wire        [(PCIE_LANE*7)-1:0] sync_fsm_rx;
 
    wire        [PCIE_LANE-1:0]     txdlysresetdone;
    wire        [PCIE_LANE-1:0]     txphaligndone;
    wire        [PCIE_LANE-1:0]     rxdlysresetdone;
    wire        [PCIE_LANE-1:0]     rxphaligndone_s;    
    
    wire                            txsyncallin;            // GTH     
    wire                            rxsyncallin;            // GTH
    
    //---------- PIPE DRP Module Output --------------------
    wire        [(PCIE_LANE*9)-1:0] drp_addr;
    wire        [PCIE_LANE-1:0]     drp_en;
    wire        [(PCIE_LANE*16)-1:0]drp_di;   
    wire        [PCIE_LANE-1:0]     drp_we;
    wire        [PCIE_LANE-1:0]     drp_done;
    wire        [(PCIE_LANE*3)-1:0] drp_fsm;

    //---------- PIPE JTAG Slave Module Output--------------
    wire	      [(PCIE_LANE*17)-1:0]jtag_sl_addr;
    wire        [PCIE_LANE-1:0]     jtag_sl_den;
    wire        [PCIE_LANE-1:0]     jtag_sl_en;
    wire        [(PCIE_LANE*16)-1:0]jtag_sl_di;
    wire        [PCIE_LANE-1:0]     jtag_sl_we;
    
    //---------- PIPE DRP MUX Output -----------------------
    wire	      [(PCIE_LANE*9)-1:0] drp_mux_addr;
    wire        [PCIE_LANE-1:0]     drp_mux_en;
    wire        [(PCIE_LANE*16)-1:0]drp_mux_di;
    wire        [PCIE_LANE-1:0]     drp_mux_we;

    //---------- PIPE EQ Module Output ---------------------
    wire        [PCIE_LANE-1:0]     eq_txeq_deemph;
    wire [(PCIE_LANE*5)-1:0] eq_txeq_precursor;
    wire        [(PCIE_LANE*7)-1:0] eq_txeq_maincursor;
    wire [(PCIE_LANE*5)-1:0] eq_txeq_postcursor;
    
    wire        [PCIE_LANE-1:0]     eq_rxeq_adapt_done;
    
    //---------- PIPE DRP Module Output --------------------
    wire        [((((PCIE_LANE-1)>>2)+1)*8)-1:0]  qdrp_addr;
    wire        [(PCIE_LANE-1)>>2:0]              qdrp_en;
    wire        [((((PCIE_LANE-1)>>2)+1)*16)-1:0] qdrp_di;   
    wire        [(PCIE_LANE-1)>>2:0]              qdrp_we;
    wire        [(PCIE_LANE-1)>>2:0]              qdrp_done;
    wire        [(PCIE_LANE-1)>>2:0]              qdrp_qpllreset;
    wire        [((((PCIE_LANE-1)>>2)+1)*6)-1:0]  qdrp_crscode;
    wire        [((((PCIE_LANE-1)>>2)+1)*9)-1:0]  qdrp_fsm;

    //---------- QPLL Wrapper Output -----------------------
    wire        [(PCIE_LANE-1)>>2:0]              qpll_qplloutclk;
    wire        [(PCIE_LANE-1)>>2:0]              qpll_qplloutrefclk;
    wire        [(PCIE_LANE-1)>>2:0]              qpll_qplllock;
    wire        [((((PCIE_LANE-1)>>2)+1)*16)-1:0] qpll_do;
    wire        [(PCIE_LANE-1)>>2:0]              qpll_rdy;

    //---------- GTX Wrapper Output ------------------------
    wire        [PCIE_LANE-1:0]     gt_txoutclk;
    wire        [PCIE_LANE-1:0]     gt_rxoutclk;
    wire        [PCIE_LANE-1:0] gt_cplllock;
    wire        [PCIE_LANE-1:0]     gt_rxcdrlock;
    wire        [PCIE_LANE-1:0]     gt_txresetdone;
    wire        [PCIE_LANE-1:0]     gt_rxresetdone;
    wire        [PCIE_LANE-1:0]     gt_eyescandataerror;
    wire        [PCIE_LANE-1:0] gt_rxpmaresetdone;
    wire        [(PCIE_LANE*8)-1:0]     gt_rxdisperr;
    wire        [(PCIE_LANE*8)-1:0]     gt_rxnotintable;
    wire        [PCIE_LANE-1:0]     gt_rxvalid;
    wire        [PCIE_LANE-1:0]     gt_phystatus;
    wire        [(PCIE_LANE*3)-1:0] gt_rxstatus;
    wire        [(PCIE_LANE*3)-1:0] gt_rxbufstatus;
    wire        [PCIE_LANE-1:0]     gt_rxelecidle;
    wire        [PCIE_LANE-1:0]     gt_txratedone;
    wire        [PCIE_LANE-1:0]     gt_rxratedone;
    wire        [(PCIE_LANE*16)-1:0]gt_do;
    wire        [PCIE_LANE-1:0]     gt_rdy;
    wire        [PCIE_LANE-1:0] gt_txphinitdone;  
    wire        [PCIE_LANE-1:0] gt_txdlysresetdone;
    wire        [PCIE_LANE-1:0] gt_txphaligndone;
    wire        [PCIE_LANE-1:0] gt_rxdlysresetdone;
    wire        [PCIE_LANE:0] gt_rxphaligndone;       // Custom width for calculation        
    wire        [PCIE_LANE-1:0]     gt_txsyncout;           // GTH  
    wire        [PCIE_LANE-1:0]     gt_txsyncdone;          // GTH                                                           
    wire        [PCIE_LANE-1:0]     gt_rxsyncout;           // GTH     
    wire        [PCIE_LANE-1:0] gt_rxsyncdone;          // GTH     
    wire        [PCIE_LANE-1:0] gt_rxcommadet;                        
    wire        [(PCIE_LANE*4)-1:0] gt_rxchariscomma;                      
    wire        [PCIE_LANE-1:0]     gt_rxbyteisaligned;                   
    wire        [PCIE_LANE-1:0]     gt_rxbyterealign; 
    wire        [ 4:0]              gt_rxchbondi [PCIE_LANE:0]; 
    wire        [(PCIE_LANE*3)-1:0] gt_rxchbondlevel;
    wire        [ 4:0]              gt_rxchbondo [PCIE_LANE:0];  
   
    wire        [PCIE_LANE-1:0]     rxchbonden;
    wire        [PCIE_LANE-1:0]     rxchbondmaster;
    wire        [PCIE_LANE-1:0]     rxchbondslave;    
    wire        [PCIE_LANE-1:0]     oobclk; 

    //---------- TX EQ -------------------------------------                                      
    localparam                      TXEQ_FS = 6'd40;        // TX equalization full swing 
    localparam                      TXEQ_LF = 6'd15;        // TX equalization low frequency

    //---------- Select JTAG Slave Type ----------------------------------------
    localparam GC_XSDB_SLAVE_TYPE = (PCIE_GT_DEVICE == "GTP") ? 16'h0400 : (PCIE_GT_DEVICE == "GTH") ? 16'h004A : 16'h0046; 

    //---------- Generate Per-Lane Signals -----------------
    genvar                          i;                      // Index for per-lane signals
    
    
    
//---------- Assignments -------------------------------------------------------
assign gt_rxchbondo[0]             = 5'd0;                  // Initialize rxchbond for lane 0 
assign gt_rxphaligndone[PCIE_LANE] = 1'd1;                  // Mot used
assign txsyncallin                 = &(gt_txphaligndone | (~user_active_lane));     
assign rxsyncallin                 = &(gt_rxphaligndone | (~user_active_lane));  

//---------- Reset Synchronizer ------------------------------------------------
always @ (posedge clk_pclk or negedge PIPE_RESET_N)
begin

    if (!PIPE_RESET_N) 
        begin
        reset_n_reg1 <= 1'd0;
        reset_n_reg2 <= 1'd0;
        end
    else
        begin
        reset_n_reg1 <= 1'd1;
        reset_n_reg2 <= reset_n_reg1;
        end   
end  


//---------- PIPE Clock Module -------------------------------------------------
generate

        begin : pipe_clock_int
model_ap2_tst_pipe_clock #
        (
        
            .PCIE_ASYNC_EN                  (PCIE_ASYNC_EN),        // PCIe async enable
            .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),        // PCIe TX buffer enable for Gen1/Gen2 only
            .PCIE_LANE                      (PCIE_LANE),            // PCIe number of lanes
            .PCIE_LINK_SPEED                (PCIE_LINK_SPEED),      // PCIe link speed 
            .PCIE_REFCLK_FREQ               (PCIE_REFCLK_FREQ),     // PCIe reference clock frequency
            .PCIE_USERCLK1_FREQ             (PCIE_USERCLK1_FREQ),   // PCIe user clock 1 frequency
            .PCIE_USERCLK2_FREQ             (PCIE_USERCLK2_FREQ),   // PCIe user clock 2 frequency
            .PCIE_OOBCLK_MODE               (PCIE_OOBCLK_MODE),     // PCIe OOB clock mode
            .PCIE_DEBUG_MODE                (PCIE_DEBUG_MODE)       // PCIe debug mode
                
        )
        model_ap2_tst_pipe_clock_i
        (
        
            //---------- Input -------------------------------------
            .CLK_CLK                        (PIPE_CLK),
            .CLK_TXOUTCLK                   (gt_txoutclk[0]),       // Reference clock from lane 0
            .CLK_RXOUTCLK_IN                (gt_rxoutclk),         
          //.CLK_RST_N                      (1'b1),                 
            .CLK_RST_N                      (PIPE_MMCM_RST_N),      // Allow system reset for error recovery             
            .CLK_PCLK_SEL                   (rate_pclk_sel),    
            .CLK_PCLK_SEL_SLAVE             (INT_PCLK_SEL_SLAVE ), 
            .CLK_GEN3                       (rate_gen3[0]),          
            
            //---------- Output ------------------------------------
            .CLK_PCLK                       (clk_pclk),
            .CLK_PCLK_SLAVE                 (INT_PCLK_OUT_SLAVE),
            .CLK_RXUSRCLK                   (clk_rxusrclk),  
            .CLK_RXOUTCLK_OUT               (clk_rxoutclk),
            .CLK_DCLK                       (clk_dclk),
            .CLK_USERCLK1                   (PIPE_USERCLK1),
            .CLK_USERCLK2                   (PIPE_USERCLK2),
            .CLK_OOBCLK                     (clk_oobclk),
            .CLK_MMCM_LOCK                  (clk_mmcm_lock)
            
        );

        assign INT_RXUSRCLK_OUT  = clk_rxusrclk;
        assign INT_RXOUTCLK_OUT  = clk_rxoutclk;
        assign INT_DCLK_OUT      = clk_dclk;
        assign INT_USERCLK1_OUT  = PIPE_USERCLK1;
        assign INT_USERCLK2_OUT  = PIPE_USERCLK2;
        assign INT_OOBCLK_OUT    = clk_oobclk;
        assign INT_MMCM_LOCK_OUT = clk_mmcm_lock;
        end 
endgenerate
   



//---------- PIPE Reset Module -------------------------------------------------
generate 

    if (PCIE_GT_DEVICE == "GTP")
        
        begin : gtp_pipe_reset

        //---------- GTP PIPE Reset Module -------------------------------------
model_ap2_tst_gtp_pipe_reset #
        (
        
            .PCIE_SIM_SPEEDUP               (PCIE_SIM_SPEEDUP),                 // PCIe sim mode
          //.PCIE_PLL_SEL                   (PCIE_PLL_SEL),                     // removed for GTP               
          //.PCIE_POWER_SAVING              (PCIE_POWER_SAVING),                // removed for GTP                                
          //.PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),                    // PCIe TX buffer enable for Gen1/Gen2 only
            .PCIE_LANE                      (PCIE_LANE)                         // PCIe number of lanes
        
        )
        model_ap2_tst_gtp_pipe_reset_i
        (
        
            //---------- Input -----------------------------
            .RST_CLK                        (clk_pclk),                 
            .RST_RXUSRCLK                   (clk_rxusrclk),
            .RST_DCLK                       (clk_dclk),
            .RST_RST_N                      (reset_n_reg2),
            .RST_DRP_DONE                   (drp_done),
            .RST_RXPMARESETDONE             (gt_rxpmaresetdone),
            .RST_PLLLOCK                    (&qpll_qplllock), 
          //.RST_QPLL_IDLE                  (qrst_idle),                        // removed for GTP  
            .RST_RATE_IDLE                  (rate_idle),
            .RST_RXCDRLOCK                  (user_rxcdrlock),
            .RST_MMCM_LOCK                  (clk_mmcm_lock),
            .RST_RESETDONE                  (user_resetdone),
            .RST_PHYSTATUS                  (gt_phystatus),
            .RST_TXSYNC_DONE                (sync_txsync_done),
            
            //---------- Output ----------------------------
            .RST_CPLLRESET                  (rst_cpllreset),                   
            .RST_CPLLPD                     (rst_cpllpd),                      
            .RST_RXUSRCLK_RESET             (rst_rxusrclk_reset),
            .RST_DCLK_RESET                 (rst_dclk_reset),
            .RST_GTRESET                    (rst_gtreset),
            .RST_DRP_START                  (rst_drp_start),
            .RST_DRP_X16                    (rst_drp_x16),
            .RST_USERRDY                    (rst_userrdy),
            .RST_TXSYNC_START               (rst_txsync_start),
            .RST_IDLE                       (rst_idle),
            .RST_FSM                        (rst_fsm)
        
        );
        
        //---------- Default ---------------------------------------------------
        assign gtp_rst_qpllreset   = rst_cpllreset;
        assign gtp_rst_qpllpd      = rst_cpllpd;
        
        end

    else 

        begin : pipe_reset

        //---------- PIPE Reset Module -----------------------------------------
model_ap2_tst_pipe_reset #
        (
        
            .PCIE_SIM_SPEEDUP               (PCIE_SIM_SPEEDUP),                 // PCIe sim mode
            .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),                   // PCIe GT Device
            .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                     // PCIe PLL select for Gen1/Gen2 only
            .PCIE_POWER_SAVING              (PCIE_POWER_SAVING),                // PCIe power saving
            .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),                    // PCIe TX buffer enable for Gen1/Gen2 only
            .PCIE_LANE                      (PCIE_LANE)                         // PCIe number of lanes
        
        )
        model_ap2_tst_pipe_reset_i
        (
        
            //---------- Input -----------------------------                    
            .RST_CLK                        (clk_pclk),                         
            .RST_RXUSRCLK                   (clk_rxusrclk),                     
            .RST_DCLK                       (clk_dclk),                         
            .RST_RST_N                      (reset_n_reg2),   
            .RST_DRP_DONE                   (drp_done),
            .RST_RXPMARESETDONE             (gt_rxpmaresetdone),                  
            .RST_CPLLLOCK                   (gt_cplllock),                      
            .RST_QPLL_IDLE                  (qrst_idle),                        
            .RST_RATE_IDLE                  (rate_idle),                        
            .RST_RXCDRLOCK                  (user_rxcdrlock),                   
            .RST_MMCM_LOCK                  (clk_mmcm_lock),                    
            .RST_RESETDONE                  (user_resetdone),                   
            .RST_PHYSTATUS                  (gt_phystatus),                     
            .RST_TXSYNC_DONE                (sync_txsync_done),                 
                                                                                
            //---------- Output ----------------------------                    
            .RST_CPLLRESET                  (rst_cpllreset),                    
            .RST_CPLLPD                     (rst_cpllpd),                       
            .RST_RXUSRCLK_RESET             (rst_rxusrclk_reset),               
            .RST_DCLK_RESET                 (rst_dclk_reset),                   
            .RST_GTRESET                    (rst_gtreset), 
            .RST_DRP_START                  (rst_drp_start),
            .RST_DRP_X16X20_MODE            (rst_drp_x16x20_mode),
            .RST_DRP_X16                    (rst_drp_x16),                     
            .RST_USERRDY                    (rst_userrdy),                      
            .RST_TXSYNC_START               (rst_txsync_start),                 
            .RST_IDLE                       (rst_idle),                         
            .RST_FSM                        (rst_fsm[4:0])                           
                                                                                
        );
       
        //---------- Default ---------------------------------------------------
        assign gtp_rst_qpllreset = 1'd0;
        assign gtp_rst_qpllpd    = 1'd0; 
       
        end
    
endgenerate



//---------- QPLL Reset Module -------------------------------------------------
generate 

    if ((PCIE_LINK_SPEED == 3) || (PCIE_PLL_SEL == "QPLL"))

        begin : qpll_reset

model_ap2_tst_qpll_reset #
        (
        
            .PCIE_PLL_SEL                   (PCIE_PLL_SEL),     // PCIe PLL select for Gen1/Gen2 only
            .PCIE_POWER_SAVING              (PCIE_POWER_SAVING),// PCIe power saving
            .PCIE_LANE                      (PCIE_LANE)         // PCIe number of lanes
            
        )
        model_ap2_tst_qpll_reset_i
        (
        
            //---------- Input ---------------------------------
            .QRST_CLK                       (clk_pclk),                 
            .QRST_RST_N                     (reset_n_reg2),
            .QRST_MMCM_LOCK                 (clk_mmcm_lock),
            .QRST_CPLLLOCK                  (gt_cplllock),
            .QRST_DRP_DONE                  (qdrp_done),
            .QRST_QPLLLOCK                  (qpll_qplllock),
            .QRST_RATE                      (PIPE_RATE),
            .QRST_QPLLRESET_IN              (rate_qpllreset),
            .QRST_QPLLPD_IN                 (rate_qpllpd),
            
            //---------- Output --------------------------------
            .QRST_OVRD                      (qrst_ovrd),
            .QRST_DRP_START                 (qrst_drp_start),
            .QRST_QPLLRESET_OUT             (qrst_qpllreset),
            .QRST_QPLLPD_OUT                (qrst_qpllpd),
            .QRST_IDLE                      (qrst_idle),
            .QRST_FSM                       (qrst_fsm)
        
        );

        end 
    
    else
     
        //---------- QPLL Reset Defaults ---------------------------------------
        begin : qpll_reset_disable
        assign qrst_ovrd      =  1'd0;
        assign qrst_drp_start =  1'd0;
        assign qrst_qpllreset =  1'd0;
        assign qrst_qpllpd    =  1'd0;
        assign qrst_idle      =  1'd0;
        assign qrst_fsm       =  1;
        end
     
endgenerate
        
assign jtag_sl_iport = {PCIE_LANE{37'd0}};

//Reference Clock for CPLLPD Fix

wire gt_cpllpdrefclk;

BUFG cpllpd_refclk_inst (.I (PIPE_CLK), .O (gt_cpllpdrefclk));

//---------- Generate PIPE Lane ------------------------------------------------
generate for (i=0; i<PCIE_LANE; i=i+1) 

    begin : pipe_lane

    //---------- PIPE User Module ----------------------------------------------
model_ap2_tst_pipe_user #
    (
    
        .PCIE_USE_MODE                  (PCIE_USE_MODE),
        .PCIE_OOBCLK_MODE               (PCIE_OOBCLK_MODE)
    
    )
    model_ap2_tst_pipe_user_i
    (
    
        //---------- Input ---------------------------------
        .USER_TXUSRCLK                  (clk_pclk),
        .USER_RXUSRCLK                  (clk_rxusrclk),
        .USER_OOBCLK_IN                 (clk_oobclk),
        .USER_RST_N                     (!rst_cpllreset),
        .USER_RXUSRCLK_RST_N            (!rst_rxusrclk_reset),
        .USER_PCLK_SEL                  (rate_pclk_sel[i]),
        .USER_RESETOVRD_START           (rate_resetovrd_start[i]),
        .USER_TXRESETDONE               (gt_txresetdone[i]),
        .USER_RXRESETDONE               (gt_rxresetdone[i]),
        .USER_TXELECIDLE                (PIPE_TXELECIDLE[i]),
        .USER_TXCOMPLIANCE              (PIPE_TXCOMPLIANCE[i]),
        .USER_RXCDRLOCK_IN              (gt_rxcdrlock[i]),
        .USER_RXVALID_IN                (gt_rxvalid[i]),
        .USER_RXSTATUS_IN               (gt_rxstatus[(3*i)+2]),
        .USER_PHYSTATUS_IN              (gt_phystatus[i]),
        .USER_RATE_DONE                 (rate_done[i]),
        .USER_RST_IDLE                  (rst_idle),
        .USER_RATE_RXSYNC               (rate_rxsync[i]),
        .USER_RATE_IDLE                 (rate_idle[i]),
        .USER_RATE_GEN3                 (rate_gen3[i]),
        .USER_RXEQ_ADAPT_DONE           (eq_rxeq_adapt_done[i]),
        
        //---------- Output --------------------------------
        .USER_OOBCLK                    (user_oobclk[i]),
        .USER_RESETOVRD                 (user_resetovrd[i]),
        .USER_TXPMARESET                (user_txpmareset[i]),                 
        .USER_RXPMARESET                (user_rxpmareset[i]),                
        .USER_RXCDRRESET                (user_rxcdrreset[i]),
        .USER_RXCDRFREQRESET            (user_rxcdrfreqreset[i]),
        .USER_RXDFELPMRESET             (user_rxdfelpmreset[i]),
        .USER_EYESCANRESET              (user_eyescanreset[i]),
        .USER_TXPCSRESET                (user_txpcsreset[i]),                   
        .USER_RXPCSRESET                (user_rxpcsreset[i]),                 
        .USER_RXBUFRESET                (user_rxbufreset[i]),
        .USER_RESETOVRD_DONE            (user_resetovrd_done[i]),
        .USER_RESETDONE                 (user_resetdone[i]),
        .USER_ACTIVE_LANE               (user_active_lane[i]),
        .USER_RXCDRLOCK_OUT             (user_rxcdrlock[i]),
        .USER_RXVALID_OUT               (PIPE_RXVALID[i]),
        .USER_PHYSTATUS_OUT             (PIPE_PHYSTATUS[i]),
        .USER_PHYSTATUS_RST             (PIPE_PHYSTATUS_RST[i]),
        .USER_GEN3_RDY                  (PIPE_GEN3_RDY[i]),
        .USER_RX_CONVERGE               (user_rx_converge[i])
    
    );
    
    
    
    //---------- GTP PIPE Rate Module ------------------------------------------
    if (PCIE_GT_DEVICE == "GTP")
    
        begin : gtp_pipe_rate
        
model_ap2_tst_gtp_pipe_rate #
       (                                                                                                           
                       
            .PCIE_SIM_SPEEDUP               (PCIE_SIM_SPEEDUP)                  // PCIe sim speedup                                                                                                        
          //.PCIE_USE_MODE                  (PCIE_USE_MODE),                    // removed for GTP                                    
          //.PCIE_PLL_SEL                   (PCIE_PLL_SEL),                     // removed for GTP               
          //.PCIE_POWER_SAVING              (PCIE_POWER_SAVING),                // removed for GTP                                
          //.PCIE_ASYNC_EN                  (PCIE_ASYNC_EN),                    // removed for GTP                               
          //.PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),                    // removed for GTP          
          //.PCIE_RXBUF_EN                  (PCIE_RXBUF_EN)                     // removed for GTP          
                                                                                                                            
        )                                                                                                           
        model_ap2_tst_gtp_pipe_rate_i
        (
    
            //---------- Input -----------------------------
            .RATE_CLK                       (clk_pclk),
            .RATE_RST_N                     (!rst_cpllreset),
          //.RATE_RST_IDLE                  (rst_idle),                         // removed for GTP
          //.RATE_ACTIVE_LANE               (user_active_lane[i]),              // removed for GTP 
            .RATE_RATE_IN                   (PIPE_RATE),   
          //.RATE_CPLLLOCK                  (gt_cplllock[i]),                   // removed for GTP
          //.RATE_QPLLLOCK                  (qpll_qplllock[i>>2])               // removed for GTP
          //.RATE_MMCM_LOCK                 (clk_mmcm_lock),                    // removed for GTP
            .RATE_DRP_DONE                  (drp_done[i]),                       
            .RATE_RXPMARESETDONE            (gt_rxpmaresetdone[i]),         
          //.RATE_TXRESETDONE               (gt_txresetdone[i]),                // removed for GTP
          //.RATE_RXRESETDONE               (gt_rxresetdone[i]),                // removed for GTP
            .RATE_TXRATEDONE                (gt_txratedone[i]),
            .RATE_RXRATEDONE                (gt_rxratedone[i]),
            .RATE_PHYSTATUS                 (gt_phystatus[i]),   
          //.RATE_RESETOVRD_DONE            (user_resetovrd_done[i]),           // removed for GTP
            .RATE_TXSYNC_DONE               (sync_txsync_done[i]),    
          //.RATE_RXSYNC_DONE               (sync_rxsync_done[i]),              // removed for GTP
                  
            //---------- Output ----------------------------
          //.RATE_CPLLPD                    (rate_cpllpd[i]),                   // removed for GTP 
          //.RATE_QPLLPD                    (rate_qpllpd[i]),                   // removed for GTP
          //.RATE_CPLLRESET                 (rate_cpllreset[i]),                // removed for GTP
          //.RATE_QPLLRESET                 (rate_qpllreset[i]),                // removed for GTP
          //.RATE_TXPMARESET                (rate_txpmareset[i]),               // removed for GTP 
          //.RATE_RXPMARESET                (rate_rxpmareset[i]),               // removed for GTP
          //.RATE_SYSCLKSEL                 (rate_sysclksel[(2*i)+1:(2*i)]),    // removed for GTP
            .RATE_DRP_START                 (rate_drp_start[i]),                
            .RATE_DRP_X16                   (rate_drp_x16[i]),
            .RATE_PCLK_SEL                  (rate_pclk_sel[i]),       
          //.RATE_GEN3                      (rate_gen3[i]),                     // removed for GTP
            .RATE_RATE_OUT                  (rate_rate[(3*i)+2:(3*i)]),      
          //.RATE_RESETOVRD_START           (rate_resetovrd_start[i]),          // removed for GTP
            .RATE_TXSYNC_START              (rate_txsync_start[i]),            
            .RATE_DONE                      (rate_done[i]),       
          //.RATE_RXSYNC_START              (rate_rxsync_start[i]),             // removed for GTP
          //.RATE_RXSYNC                    (rate_rxsync[i]),                   // removed for GTP
            .RATE_IDLE                      (rate_idle[i]),                     
            .RATE_FSM                       (rate_fsm[(5*i)+4:(5*i)])       
        );
    
        //---------- Default for GTP -----------------------
        assign rate_cpllpd[i]                = 1'd0;
        assign rate_qpllpd[i]                = 1'd0;
        assign rate_cpllreset[i]             = 1'd0;
        assign rate_qpllreset[i]             = 1'd0;
        assign rate_txpmareset[i]            = 1'd0;
        assign rate_rxpmareset[i]            = 1'd0;
        assign rate_sysclksel[(2*i)+1:(2*i)] = 2'b0;
        assign rate_gen3[i]                  = 1'd0;
        assign rate_resetovrd_start[i]       = 1'd0;
        assign rate_rxsync_start[i]          = 1'd0;
        assign rate_rxsync[i]                = 1'd0; 
        
        end 
    
    else
    
        begin : pipe_rate
    
        //---------- PIPE Rate Module ----------------------------------------------                                     
model_ap2_tst_pipe_rate #
        (
        
            .PCIE_SIM_SPEEDUP               (PCIE_SIM_SPEEDUP), // PCIe sim speedup 
            .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),   // PCIe GT device
            .PCIE_USE_MODE                  (PCIE_USE_MODE),    // PCIe use mode
            .PCIE_PLL_SEL                   (PCIE_PLL_SEL),     // PCIe PLL select for Gen1/Gen2 only
            .PCIE_POWER_SAVING              (PCIE_POWER_SAVING),// PCIe power saving
            .PCIE_ASYNC_EN                  (PCIE_ASYNC_EN),    // PCIe async enable
            .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),    // PCIe TX buffer enable for Gen1/Gen2 only
            .PCIE_RXBUF_EN                  (PCIE_RXBUF_EN)     // PCIe RX buffer enable for Gen3      only
            
        )
        model_ap2_tst_pipe_rate_i
        (
        
            //---------- Input ---------------------------------                                
            .RATE_CLK                       (clk_pclk),                                         
            .RATE_RST_N                     (!rst_cpllreset),                                   
            .RATE_RST_IDLE                  (rst_idle),                                         
            .RATE_ACTIVE_LANE               (user_active_lane[i]),                              
            .RATE_RATE_IN                   (PIPE_RATE),                                        
            .RATE_CPLLLOCK                  (gt_cplllock[i]),                                   
            .RATE_QPLLLOCK                  (qpll_qplllock[i>>2]),                              
            .RATE_MMCM_LOCK                 (clk_mmcm_lock),                                    
            .RATE_DRP_DONE                  (drp_done[i]),      
            .RATE_RXPMARESETDONE            (gt_rxpmaresetdone[i]),                                
            .RATE_TXRESETDONE               (gt_txresetdone[i]),                                
            .RATE_RXRESETDONE               (gt_rxresetdone[i]),                                
            .RATE_TXRATEDONE                (gt_txratedone[i]),                                 
            .RATE_RXRATEDONE                (gt_rxratedone[i]),                                 
            .RATE_PHYSTATUS                 (gt_phystatus[i]),                                  
            .RATE_RESETOVRD_DONE            (user_resetovrd_done[i]),                           
            .RATE_TXSYNC_DONE               (sync_txsync_done[i]),        		                  
            .RATE_RXSYNC_DONE               (sync_rxsync_done[i]),	                            
                                                                                                
            //---------- Output --------------------------------                                
            .RATE_CPLLPD                    (rate_cpllpd[i]),                                   
            .RATE_QPLLPD                    (rate_qpllpd[i]),                                   
            .RATE_CPLLRESET                 (rate_cpllreset[i]),                                
            .RATE_QPLLRESET                 (rate_qpllreset[i]),                                
            .RATE_TXPMARESET                (rate_txpmareset[i]),                               
            .RATE_RXPMARESET                (rate_rxpmareset[i]),                               
            .RATE_SYSCLKSEL                 (rate_sysclksel[(2*i)+1:(2*i)]),                    
            .RATE_DRP_START                 (rate_drp_start[i]),  
            .RATE_DRP_X16X20_MODE           (rate_drp_x16x20_mode[i]),      
            .RATE_DRP_X16                   (rate_drp_x16[i]),                        
            .RATE_PCLK_SEL                  (rate_pclk_sel[i]),                                 
            .RATE_GEN3                      (rate_gen3[i]),                                     
            .RATE_RATE_OUT                  (rate_rate[(3*i)+2:(3*i)]),                         
            .RATE_RESETOVRD_START           (rate_resetovrd_start[i]),
            .RATE_TXSYNC_START              (rate_txsync_start[i]),
            .RATE_DONE                      (rate_done[i]),
            .RATE_RXSYNC_START              (rate_rxsync_start[i]),
            .RATE_RXSYNC                    (rate_rxsync[i]),
            .RATE_IDLE                      (rate_idle[i]),
            .RATE_FSM                       (rate_fsm[(5*i)+4:(5*i)])
            
        );    
        
        end
    
    
    
    //---------- PIPE Sync Module ----------------------------------------------
model_ap2_tst_pipe_sync #
    (
    
        .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),   // PCIe GT Device
        .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),    // PCIe TX buffer enable for Gen1/Gen2 only
        .PCIE_RXBUF_EN                  (PCIE_RXBUF_EN),    // PCIe RX buffer enable for Gen3      only
        .PCIE_TXSYNC_MODE               (PCIE_TXSYNC_MODE), // PCIe TX sync mode
        .PCIE_RXSYNC_MODE               (PCIE_RXSYNC_MODE), // PCIe RX sync mode
        .PCIE_LANE                      (PCIE_LANE),        // PCIe lane
        .PCIE_LINK_SPEED                (PCIE_LINK_SPEED)   // PCIe link speed
    
    )
    model_ap2_tst_pipe_sync_i 
    (
    
        //---------- Input ---------------------------------
        .SYNC_CLK                       (clk_pclk),
        .SYNC_RST_N                     (!rst_cpllreset),
        .SYNC_SLAVE                     (i > 0),
        .SYNC_GEN3                      (rate_gen3[i]),
        .SYNC_RATE_IDLE                 (rate_idle[i]),
        .SYNC_MMCM_LOCK                 (clk_mmcm_lock),
        .SYNC_RXELECIDLE                (gt_rxelecidle[i]),
        .SYNC_RXCDRLOCK                 (user_rxcdrlock[i]),
        .SYNC_ACTIVE_LANE               (user_active_lane[i]),
        
        .SYNC_TXSYNC_START              (rate_txsync_start[i] || rst_txsync_start),
        .SYNC_TXPHINITDONE              (&(gt_txphinitdone | (~user_active_lane))),     
        .SYNC_TXDLYSRESETDONE           (txdlysresetdone[i]),                 
        .SYNC_TXPHALIGNDONE             (txphaligndone[i]),  
        .SYNC_TXSYNCDONE                (gt_txsyncdone[i]), // GTH
        
        .SYNC_RXSYNC_START              (rate_rxsync_start[i]),
        .SYNC_RXDLYSRESETDONE           (rxdlysresetdone[i]),
        .SYNC_RXPHALIGNDONE_M           (gt_rxphaligndone[0]),
        .SYNC_RXPHALIGNDONE_S           (rxphaligndone_s[i]),
        .SYNC_RXSYNC_DONEM_IN           (sync_rxsync_donem[0]),   
        .SYNC_RXSYNCDONE                (gt_rxsyncdone[i]), // GTH
    
        //---------- Output --------------------------------
        .SYNC_TXPHDLYRESET              (sync_txphdlyreset[i]),
        .SYNC_TXPHALIGN                 (sync_txphalign[i]),           
        .SYNC_TXPHALIGNEN               (sync_txphalignen[i]),        
        .SYNC_TXPHINIT                  (sync_txphinit[i]),    
        .SYNC_TXDLYBYPASS               (sync_txdlybypass[i]),                   
        .SYNC_TXDLYSRESET               (sync_txdlysreset[i]),
        .SYNC_TXDLYEN                   (sync_txdlyen[i]), 
        .SYNC_TXSYNC_DONE               (sync_txsync_done[i]),
        .SYNC_FSM_TX                    (sync_fsm_tx[(6*i)+5:(6*i)]),
        
        .SYNC_RXPHALIGN                 (sync_rxphalign[i]),
        .SYNC_RXPHALIGNEN               (sync_rxphalignen[i]),
        .SYNC_RXDLYBYPASS               (sync_rxdlybypass[i]),          
        .SYNC_RXDLYSRESET               (sync_rxdlysreset[i]),
        .SYNC_RXDLYEN                   (sync_rxdlyen[i]),
        .SYNC_RXDDIEN                   (sync_rxddien[i]),
        .SYNC_RXSYNC_DONEM_OUT          (sync_rxsync_donem[i]),
        .SYNC_RXSYNC_DONE               (sync_rxsync_done[i]),
        .SYNC_FSM_RX                    (sync_fsm_rx[(7*i)+6:(7*i)])
        
    );
    
    //---------- PIPE Sync Assignments -----------------------------------------
    assign txdlysresetdone[i] = (PCIE_TXSYNC_MODE == 1) ? gt_txdlysresetdone[i] : &gt_txdlysresetdone;
    assign txphaligndone[i]   = (PCIE_TXSYNC_MODE == 1) ? gt_txphaligndone[i]   : &(gt_txphaligndone | (~user_active_lane));
    assign rxdlysresetdone[i] = (PCIE_RXSYNC_MODE == 1) ? gt_rxdlysresetdone[i] : &gt_rxdlysresetdone;
    assign rxphaligndone_s[i] = (PCIE_LANE == 1)        ? 1'd0                  : &gt_rxphaligndone[PCIE_LANE:1];
    
    
    //---------- GTP PIPE DRP Module -------------------------------------------
    if (PCIE_GT_DEVICE == "GTP")
    
        begin : gtp_pipe_drp
       
        //---------- GTP PIPE DRP Module ---------------------------------------
model_ap2_tst_gtp_pipe_drp 
        model_ap2_tst_gtp_pipe_drp_i
        (
            
            //---------- Input ---------------------------------
            .DRP_CLK                        (clk_dclk),
            .DRP_RST_N                      (!rst_dclk_reset),
            .DRP_X16                        (rst_drp_x16 || rate_drp_x16[i]),
            .DRP_START                      (rst_drp_start || rate_drp_start[i]),                      
            .DRP_DO                         (gt_do[(16*i)+15:(16*i)]),
            .DRP_RDY                        (gt_rdy[i]),
            
            //---------- Output --------------------------------
            .DRP_ADDR                       (drp_addr[(9*i)+8:(9*i)]),
            .DRP_EN                         (drp_en[i]),  
            .DRP_DI                         (drp_di[(16*i)+15:(16*i)]),   
            .DRP_WE                         (drp_we[i]),
            .DRP_DONE                       (drp_done[i]),
            .DRP_FSM                        (drp_fsm[(3*i)+2:(3*i)])
            
        );
        
        end
       
    else
    
        begin : pipe_drp 
        
        //---------- PIPE DRP Module -------------------------------------------
model_ap2_tst_pipe_drp #
        (
        
            .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),                   // PCIe GT device
            .PCIE_USE_MODE                  (PCIE_USE_MODE),                    // PCIe use mode
            .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                     // PCIe PLL select for Gen1/Gen2 only
            .PCIE_AUX_CDR_GEN3_EN           (PCIE_AUX_CDR_GEN3_EN),             // PCIe AUX CDR Gen3 enable
            .PCIE_ASYNC_EN                  (PCIE_ASYNC_EN),                    // PCIe async enable
            .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),                    // PCIe TX buffer enable for Gen1/Gen2 only
            .PCIE_RXBUF_EN                  (PCIE_RXBUF_EN),                    // PCIe RX buffer enable for Gen3      only
            .PCIE_TXSYNC_MODE               (PCIE_TXSYNC_MODE),                 // PCIe TX sync mode
            .PCIE_RXSYNC_MODE               (PCIE_RXSYNC_MODE)                  // PCIe RX sync mode
        
        )
        model_ap2_tst_pipe_drp_i
        (
            
            //---------- Input ---------------------------------
            .DRP_CLK                        (clk_dclk),
            .DRP_RST_N                      (!rst_dclk_reset),
            .DRP_GTXRESET                   (rst_gtreset),
            .DRP_RATE                       (PIPE_RATE),
            .DRP_X16X20_MODE                (rst_drp_x16x20_mode || rate_drp_x16x20_mode[i]),
            .DRP_X16                        (rst_drp_x16         || rate_drp_x16[i]),
            .DRP_START                      (rst_drp_start || rate_drp_start[i]),                      
            .DRP_DO                         (gt_do[(16*i)+15:(16*i)]),
            .DRP_RDY                        (gt_rdy[i]),
            
            //---------- Output --------------------------------
            .DRP_ADDR                       (drp_addr[(9*i)+8:(9*i)]),
            .DRP_EN                         (drp_en[i]),  
            .DRP_DI                         (drp_di[(16*i)+15:(16*i)]),   
            .DRP_WE                         (drp_we[i]),
            .DRP_DONE                       (drp_done[i]),
            .DRP_FSM                        (drp_fsm[(3*i)+2:(3*i)])
            
        );
        
        end

    
         assign jtag_sl_oport[((i+1)*17)-1 : (i*17)] = 17'd0;
         assign jtag_sl_addr[(17*i)+16:(17*i)]       = 17'd0;   
         assign jtag_sl_den[i]                       =  1'd0;
         assign jtag_sl_di[(16*i)+15:(16*i)]         = 16'd0;
         assign jtag_sl_we[i]                        =  1'd0;

    //---------- Generate DRP MUX ----------------------------------------------
    assign PIPE_JTAG_RDY[i] = (drp_fsm[(3*i)+2:(3*i)] == 3'b000);
    assign jtag_sl_en[i]	  = (jtag_sl_addr[(17*i)+16:(17*i)+9] == 8'd0) ? jtag_sl_den[i] : 1'd0;

    // Channel DRP
    assign drp_mux_en[i]                = (PIPE_JTAG_RDY[i] && EXT_CH_GT_DRP) ? EXT_CH_GT_DRPEN[i] : drp_en[i];
    assign drp_mux_di[(16*i)+15:(16*i)] = (PIPE_JTAG_RDY[i] && EXT_CH_GT_DRP) ? EXT_CH_GT_DRPDI[(16*i)+15:(16*i)] : drp_di[(16*i)+15:(16*i)];
    assign drp_mux_addr[(9*i)+8:(9*i)]  = (PIPE_JTAG_RDY[i] && EXT_CH_GT_DRP) ? EXT_CH_GT_DRPADDR[(9*i)+8:(9*i)] : drp_addr[(9*i)+8:(9*i)];
    assign drp_mux_we[i]                = (PIPE_JTAG_RDY[i] && EXT_CH_GT_DRP) ? EXT_CH_GT_DRPWE[i]  : drp_we[i];

    //---------- Generate PIPE EQ ----------------------------------------------
    if (PCIE_LINK_SPEED == 3) 
    
        begin : pipe_eq
    
        //---------- PIPE EQ Module --------------------------------------------
model_ap2_tst_pipe_eq #
        (
            .PCIE_SIM_MODE                  (PCIE_SIM_MODE),                    // PCIe sim mode
            .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),
            .PCIE_RXEQ_MODE_GEN3            (PCIE_RXEQ_MODE_GEN3)               // PCIe RX equalization mode
        )
        model_ap2_tst_pipe_eq_i
        (
        
            //---------- Input -----------------------------
            .EQ_CLK                         (clk_pclk),
            .EQ_RST_N                       (!rst_cpllreset),
            .EQ_GEN3                        (rate_gen3[i]),
            
            .EQ_TXEQ_CONTROL                (PIPE_TXEQ_CONTROL[(2*i)+1:(2*i)]),    
            .EQ_TXEQ_PRESET                 (PIPE_TXEQ_PRESET[(4*i)+3:(4*i)]),
            .EQ_TXEQ_PRESET_DEFAULT         (PIPE_TXEQ_PRESET_DEFAULT[(4*i)+3:(4*i)]),
            .EQ_TXEQ_DEEMPH_IN              (PIPE_TXEQ_DEEMPH[(6*i)+5:(6*i)]),  // renamed
                                           
            .EQ_RXEQ_CONTROL                (PIPE_RXEQ_CONTROL[(2*i)+1:(2*i)]),  
            .EQ_RXEQ_PRESET                 (PIPE_RXEQ_PRESET[(3*i)+2:(3*i)]),
            .EQ_RXEQ_LFFS                   (PIPE_RXEQ_LFFS[(6*i)+5:(6*i)]),  
            .EQ_RXEQ_TXPRESET               (PIPE_RXEQ_TXPRESET[(4*i)+3:(4*i)]),
            .EQ_RXEQ_USER_EN                (PIPE_RXEQ_USER_EN[i]),          
            .EQ_RXEQ_USER_TXCOEFF           (PIPE_RXEQ_USER_TXCOEFF[(18*i)+17:(18*i)]),     
            .EQ_RXEQ_USER_MODE              (PIPE_RXEQ_USER_MODE[i]),        
            
            //---------- Output ----------------------------
            .EQ_TXEQ_DEEMPH                 (eq_txeq_deemph[i]),
            .EQ_TXEQ_PRECURSOR              (eq_txeq_precursor[(5*i)+4:(5*i)]),
            .EQ_TXEQ_MAINCURSOR             (eq_txeq_maincursor[(7*i)+6:(7*i)]),
            .EQ_TXEQ_POSTCURSOR             (eq_txeq_postcursor[(5*i)+4:(5*i)]),
            .EQ_TXEQ_DEEMPH_OUT             (PIPE_TXEQ_COEFF[(18*i)+17:(18*i)]),// renamed
            .EQ_TXEQ_DONE                   (PIPE_TXEQ_DONE[i]),
            .EQ_TXEQ_FSM                    (PIPE_TXEQ_FSM[(6*i)+5:(6*i)]),
            
            .EQ_RXEQ_NEW_TXCOEFF            (PIPE_RXEQ_NEW_TXCOEFF[(18*i)+17:(18*i)]), 
            .EQ_RXEQ_LFFS_SEL               (PIPE_RXEQ_LFFS_SEL[i]),
            .EQ_RXEQ_ADAPT_DONE             (eq_rxeq_adapt_done[i]),
            .EQ_RXEQ_DONE                   (PIPE_RXEQ_DONE[i]),
            .EQ_RXEQ_FSM                    (PIPE_RXEQ_FSM[(6*i)+5:(6*i)])
        
        );
    
        end 
        
    else
    
        //---------- PIPE EQ Defaults ------------------------------------------
        begin : pipe_eq_disable                      
        assign eq_txeq_deemph[i]                       =  1'd0;
        assign eq_txeq_precursor[(5*i)+4:(5*i)]        =  5'h00;
        assign eq_txeq_maincursor[(7*i)+6:(7*i)]       =  7'h00;
        assign eq_txeq_postcursor[(5*i)+4:(5*i)]       =  5'h00;
        assign eq_rxeq_adapt_done[i]                   =  1'd0;
        assign PIPE_TXEQ_COEFF[(18*i)+17:(18*i)]       = 18'd0;
        assign PIPE_TXEQ_DONE[i]                       =  1'd0;
        assign PIPE_TXEQ_FSM[(6*i)+5:(6*i)]            =  6'd0;
        
        assign PIPE_RXEQ_NEW_TXCOEFF[(18*i)+17:(18*i)] = 18'd0;
        assign PIPE_RXEQ_LFFS_SEL[i]                   =  1'd0;
        assign PIPE_RXEQ_ADAPT_DONE[i]                 =  1'd0;   
        assign PIPE_RXEQ_DONE[i]                       =  1'd0;                                     
        assign PIPE_RXEQ_FSM[(6*i)+5:(6*i)]            =  6'd0;   
        end

    //---------- Generate PIPE Common Per Quad for Gen3 ------------------------
    if ((i%4)==0)

        begin : pipe_quad

        //---------- Generate QPLL Powerdown and Reset -------------------------
        assign qpllpd          = (PCIE_GT_DEVICE == "GTP") ? gtp_rst_qpllpd    : qrst_qpllpd;
        assign qpllreset[i>>2] = (PCIE_GT_DEVICE == "GTP") ? gtp_rst_qpllreset : (qrst_qpllreset || qdrp_qpllreset[i>>2]);

        if ((PCIE_LINK_SPEED == 3) || (PCIE_PLL_SEL == "QPLL") || (PCIE_GT_DEVICE == "GTP"))

           begin : gt_common_enabled

           if (PCIE_EXT_GT_COMMON == "FALSE")

           begin : gt_common_int

    //---------- GT COMMON INTERNAL Module ---------------------------------------
model_ap2_tst_gt_common #
            (

                .PCIE_SIM_MODE                  (PCIE_SIM_MODE),                // PCIe sim mode
                .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),               // PCIe GT device
                .PCIE_USE_MODE                  (PCIE_USE_MODE),                // PCIe use mode
                .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                 // PCIe PLL select for Gen1/Gen2 only
                .PCIE_REFCLK_FREQ               (PCIE_REFCLK_FREQ)              // PCIe reference clock frequency

            )
            model_ap2_tst_gt_common_i
            (

                //---------- Input -------------------------
                .CPLLPDREFCLK                        (gt_cpllpdrefclk),
                .PIPE_CLK                            (PIPE_CLK),
                .QPLL_QPLLPD                         (qpllpd),
                .QPLL_QPLLRESET                      (qpllreset[i>>2]),
                .QPLL_DRP_CLK                        (clk_dclk),
                .QPLL_DRP_RST_N                      (rst_dclk_reset),
                .QPLL_DRP_OVRD                       (qrst_ovrd),
                .QPLL_DRP_GEN3                       (&rate_gen3),
                .QPLL_DRP_START                      (qrst_drp_start),

                .QPLL_DRP_CRSCODE                    (qdrp_crscode[(6*(i>>2))+5:(6*(i>>2))]),
                .QPLL_DRP_FSM                        (qdrp_fsm[(9*(i>>2))+8:(9*(i>>2))]),
                .QPLL_DRP_DONE                       (qdrp_done[i>>2]),
                .QPLL_DRP_RESET                      (qdrp_qpllreset[i>>2]),
                .QPLL_QPLLOUTCLK                     (qpll_qplloutclk[i>>2]),
                .QPLL_QPLLOUTREFCLK                  (qpll_qplloutrefclk[i>>2]),
                .QPLL_QPLLLOCK                       (qpll_qplllock[i>>2])
            );
              assign QPLL_QPLLPD                           =  1'b0;
              assign QPLL_QPLLRESET[i>>2]                  =  1'b0;              
              assign QPLL_DRP_CLK                          =  1'b0;
              assign QPLL_DRP_RST_N                        =  1'b0;
              assign QPLL_DRP_OVRD                         =  1'b0;
              assign QPLL_DRP_GEN3                         =  1'b0;
              assign QPLL_DRP_START                        =  1'b0;
              assign INT_QPLLLOCK_OUT[i>>2]                =  qpll_qplllock[i>>2] ;
              assign INT_QPLLOUTREFCLK_OUT[i>>2]           =  qpll_qplloutrefclk[i>>2];
              assign INT_QPLLOUTCLK_OUT[i>>2]              =  qpll_qplloutclk[i>>2];
            end
         else
            begin   : gt_common_ext
              assign qdrp_done[i>>2]                       =  QPLL_DRP_DONE[i>>2];
              assign qdrp_qpllreset[i>>2]                  =  QPLL_DRP_RESET[i>>2];
              assign qdrp_crscode[(6*(i>>2))+5:(6*(i>>2))] =  QPLL_DRP_CRSCODE[(6*(i>>2))+5:(6*(i>>2))];
              assign qdrp_fsm[(9*(i>>2))+8:(9*(i>>2))]     =  QPLL_DRP_FSM[(9*(i>>2))+8:(9*(i>>2))];
              assign qpll_qplloutclk[i>>2]                 =  QPLL_QPLLOUTCLK[i>>2];
              assign qpll_qplloutrefclk[i>>2]              =  QPLL_QPLLOUTREFCLK[i>>2];
              assign qpll_qplllock[i>>2]                   =  QPLL_QPLLLOCK[i>>2];
              assign QPLL_QPLLPD                           =  qpllpd;
              assign QPLL_QPLLRESET[i>>2]                  =  qpllreset[i>>2];              
              assign QPLL_DRP_CLK                          =  clk_dclk;
              assign QPLL_DRP_RST_N                        =  rst_dclk_reset;
              assign QPLL_DRP_OVRD                         =  qrst_ovrd;
              assign QPLL_DRP_GEN3                         =  &rate_gen3;
              assign QPLL_DRP_START                        =  qrst_drp_start;
              assign INT_QPLLLOCK_OUT[i>>2]                =  1'b0;
              assign INT_QPLLOUTCLK_OUT[i>>2]              =  1'b0;
              assign INT_QPLLOUTREFCLK_OUT[i>>2]           =  1'b0;
            end
         end
       else

            //---------- PIPE Common Defaults ----------------------------------
            begin : gt_common_disabled
            assign qdrp_done[i>>2]                       =  1'd0;
            assign qdrp_crscode[(6*(i>>2))+5:(6*(i>>2))] =  6'd0;
            assign qdrp_fsm[(9*(i>>2))+8:(9*(i>>2))]     =  9'd0;
            assign qpll_qplloutclk[i>>2]                 =  1'd0;
            assign qpll_qplloutrefclk[i>>2]              =  1'd0;
            assign qpll_qplllock[i>>2]                   =  1'd0;
            assign QPLL_QPLLPD                           =  1'b0;
            assign QPLL_QPLLRESET[i>>2]                  =  1'b0;              
            assign QPLL_DRP_CLK                          =  1'b0;
            assign QPLL_DRP_RST_N                        =  1'b0;
            assign QPLL_DRP_OVRD                         =  1'b0;
            assign QPLL_DRP_GEN3                         =  1'b0;
            assign QPLL_DRP_START                        =  1'b0;
            assign INT_QPLLLOCK_OUT[i>>2]                =  1'b0;
            assign INT_QPLLOUTCLK_OUT[i>>2]              =  1'b0;
            assign INT_QPLLOUTREFCLK_OUT[i>>2]           =  1'b0;
            end
     end

    //---------- GT Wrapper ----------------------------------------------------
    assign gt_txpmareset_i[i] = (user_txpmareset[i] || rate_txpmareset[i]);
    assign gt_rxpmareset_i[i] = (user_rxpmareset[i] || rate_rxpmareset[i]);

model_ap2_tst_gt_wrapper #
    (
    
        .PCIE_SIM_MODE                  (PCIE_SIM_MODE),                        // PCIe sim mode
        .PCIE_SIM_SPEEDUP               (PCIE_SIM_SPEEDUP),                     // PCIe sim speedup
        .PCIE_SIM_TX_EIDLE_DRIVE_LEVEL  (PCIE_SIM_TX_EIDLE_DRIVE_LEVEL),        // PCIe sim TX electrical idle drive level 
        .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),                       // PCIe GT device
        .PCIE_USE_MODE                  (PCIE_USE_MODE),                        // PCIe use mode
        .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                         // PCIe PLL select for Gen1/Gen2 only
        .PCIE_LPM_DFE                   (PCIE_LPM_DFE),                         // PCIe LPM or DFE mode for Gen1/Gen2 only
        .PCIE_LPM_DFE_GEN3              (PCIE_LPM_DFE_GEN3),                    // PCIe LPM or DFE mode for Gen3      only
        .PCIE_ASYNC_EN                  (PCIE_ASYNC_EN),                        // PCIe async enable
        .PCIE_TXBUF_EN                  (PCIE_TXBUF_EN),                        // PCIe TX buffer enable for Gen1/Gen2 only
        .PCIE_TXSYNC_MODE               (PCIE_TXSYNC_MODE),                     // PCIe TX sync mode
        .PCIE_RXSYNC_MODE               (PCIE_RXSYNC_MODE),                     // PCIe RX sync mode
        .PCIE_CHAN_BOND                 (PCIE_CHAN_BOND),                       // PCIe Channel bonding mode
        .PCIE_CHAN_BOND_EN              (PCIE_CHAN_BOND_EN),                    // PCIe Channel bonding enable for Gen1/Gen2 only
        .PCIE_LANE                      (PCIE_LANE),                            // PCIe number of lane
        .PCIE_REFCLK_FREQ               (PCIE_REFCLK_FREQ),                     // PCIe reference clock frequency
        .PCIE_TX_EIDLE_ASSERT_DELAY     (PCIE_TX_EIDLE_ASSERT_DELAY),           // PCIe TX electrical idle assert delay
        .PCIE_OOBCLK_MODE               (PCIE_OOBCLK_MODE),                     // PCIe OOB clock mode
        .TX_MARGIN_FULL_0               (TX_MARGIN_FULL_0),                      
        .TX_MARGIN_FULL_1               (TX_MARGIN_FULL_1),   
        .TX_MARGIN_FULL_2               (TX_MARGIN_FULL_2),
        .TX_MARGIN_FULL_3               (TX_MARGIN_FULL_3),
        .TX_MARGIN_FULL_4               (TX_MARGIN_FULL_4),
        .TX_MARGIN_LOW_0                (TX_MARGIN_LOW_0), 
        .TX_MARGIN_LOW_1                (TX_MARGIN_LOW_1), 
        .TX_MARGIN_LOW_2                (TX_MARGIN_LOW_2),
        .TX_MARGIN_LOW_3                (TX_MARGIN_LOW_3),
        .TX_MARGIN_LOW_4                (TX_MARGIN_LOW_4),

        .PCIE_DEBUG_MODE                (PCIE_DEBUG_MODE)                       // PCIe debug mode
    )
    model_ap2_tst_gt_wrapper_i
    (
    
        //---------- GT User Ports -------------------------
        .GT_MASTER                      (i == 0),
        .GT_GEN3                        (rate_gen3[i]),   
        .GT_RX_CONVERGE                 (&user_rx_converge),     
    
        //---------- GT Clock Ports ------------------------
        .GT_GTREFCLK0                   (PIPE_CLK),
        .GT_QPLLCLK                     (qpll_qplloutclk[i>>2]),
        .GT_QPLLREFCLK                  (qpll_qplloutrefclk[i>>2]),
        .GT_TXUSRCLK                    (clk_pclk),
        .GT_RXUSRCLK                    (clk_rxusrclk), 
        .GT_TXUSRCLK2                   (clk_pclk),
        .GT_RXUSRCLK2                   (clk_rxusrclk), 
        .GT_OOBCLK                      (oobclk[i]),
        .GT_TXSYSCLKSEL                 (rate_sysclksel[(2*i)+1:(2*i)]),
        .GT_RXSYSCLKSEL                 (rate_sysclksel[(2*i)+1:(2*i)]),
        .GT_CPLLPDREFCLK                (gt_cpllpdrefclk),
                                
        .GT_TXOUTCLK                    (gt_txoutclk[i]),
        .GT_RXOUTCLK                    (gt_rxoutclk[i]),
        .GT_CPLLLOCK                    (gt_cplllock[i]),  
        .GT_RXCDRLOCK                   (gt_rxcdrlock[i]),
        
        //---------- GT Reset Ports ------------------------
        .GT_CPLLPD                      (rst_cpllpd    || rate_cpllpd[i]),
        .GT_CPLLRESET                   (rst_cpllreset || rate_cpllreset[i]),
        .GT_TXUSERRDY                   (rst_userrdy),
        .GT_RXUSERRDY                   (rst_userrdy),
        .GT_RESETOVRD                   (user_resetovrd[i]),
        .GT_GTTXRESET                   (rst_gtreset),
        .GT_GTRXRESET                   (rst_gtreset),
        .GT_TXPMARESET                  (gt_txpmareset_i[i]), // (user_txpmareset[i] || rate_txpmareset[i]),                 
        .GT_RXPMARESET                  (gt_rxpmareset_i[i]), // (user_rxpmareset[i] || rate_rxpmareset[i]),                
        .GT_RXCDRRESET                  (user_rxcdrreset[i]),
        .GT_RXCDRFREQRESET              (user_rxcdrfreqreset[i]),
        .GT_RXDFELPMRESET               (user_rxdfelpmreset[i]),
        .GT_EYESCANRESET                (user_eyescanreset[i]),
        .GT_TXPCSRESET                  (user_txpcsreset[i]),                   
        .GT_RXPCSRESET                  (user_rxpcsreset[i]),                 
        .GT_RXBUFRESET                  (user_rxbufreset[i]),
                                    
        .GT_EYESCANDATAERROR            (gt_eyescandataerror[i]),
        .GT_TXRESETDONE                 (gt_txresetdone[i]),
        .GT_RXRESETDONE                 (gt_rxresetdone[i]),
        .GT_RXPMARESETDONE              (gt_rxpmaresetdone[i]),
        
        //---------- GT TX Data Ports ----------------------
        .GT_TXDATA                      (PIPE_TXDATA[(32*i)+31:(32*i)]),
        .GT_TXDATAK                     (PIPE_TXDATAK[(4*i)+3:(4*i)]),
        
        .GT_TXP                         (PIPE_TXP[i]),
        .GT_TXN                         (PIPE_TXN[i]),
        
        //---------- GT RX Data Ports ----------------------
        .GT_RXP                         (PIPE_RXP[i]),
        .GT_RXN                         (PIPE_RXN[i]),
        
        .GT_RXDATA                      (PIPE_RXDATA[(32*i)+31:(32*i)]),
        .GT_RXDATAK                     (PIPE_RXDATAK[(4*i)+3:(4*i)]),
        
        //---------- GT Command Ports ----------------------
        .GT_TXDETECTRX                  (PIPE_TXDETECTRX),
        .GT_TXELECIDLE                  (PIPE_TXELECIDLE[i]), 
        .GT_TXCOMPLIANCE                (PIPE_TXCOMPLIANCE[i]),
        .GT_RXPOLARITY                  (PIPE_RXPOLARITY[i]),
        .GT_TXPOWERDOWN                 (PIPE_POWERDOWN[(2*i)+1:(2*i)]),
        .GT_RXPOWERDOWN                 (PIPE_POWERDOWN[(2*i)+1:(2*i)]),
        .GT_TXRATE                      (rate_rate[(3*i)+2:(3*i)]),
        .GT_RXRATE                      (rate_rate[(3*i)+2:(3*i)]),        
            
        //---------- GT Electrical Command Ports -----------
        .GT_TXMARGIN                    (PIPE_TXMARGIN),
        .GT_TXSWING                     (PIPE_TXSWING),
        .GT_TXDEEMPH                    (PIPE_TXDEEMPH[i]),  
        .GT_TXPRECURSOR                 (eq_txeq_precursor[(5*i)+4:(5*i)]),
        .GT_TXMAINCURSOR                (eq_txeq_maincursor[(7*i)+6:(7*i)]),
        .GT_TXPOSTCURSOR                (eq_txeq_postcursor[(5*i)+4:(5*i)]),
    
        //---------- GT Status Ports -----------------------
        .GT_RXVALID                     (gt_rxvalid[i]),
        .GT_PHYSTATUS                   (gt_phystatus[i]),
        .GT_RXELECIDLE                  (gt_rxelecidle[i]),
        .GT_RXSTATUS                    (gt_rxstatus[(3*i)+2:(3*i)]),
        .GT_RXBUFSTATUS                 (gt_rxbufstatus[(3*i)+2:(3*i)]),
        .GT_TXRATEDONE                  (gt_txratedone[i]),
        .GT_RXRATEDONE                  (gt_rxratedone[i]),
        .GT_RXDISPERR                   (gt_rxdisperr[(8*i)+7:(8*i)]),  
        .GT_RXNOTINTABLE                (gt_rxnotintable[(8*i)+7:(8*i)]),
    
        //---------- GT DRP Ports --------------------------
        .GT_DRPCLK                      (clk_dclk),
        .GT_DRPADDR                     (drp_mux_addr[(9*i)+8:(9*i)]),
        .GT_DRPEN                       (drp_mux_en[i]),
        .GT_DRPDI                       (drp_mux_di[(16*i)+15:(16*i)]),
        .GT_DRPWE                       (drp_mux_we[i]),
                                     
        .GT_DRPDO                       (gt_do[(16*i)+15:(16*i)]),
        .GT_DRPRDY                      (gt_rdy[i]),
        
        //---------- GT TX Sync Ports ----------------------
        .GT_TXPHALIGN                   (sync_txphalign[i]),    
        .GT_TXPHALIGNEN                 (sync_txphalignen[i]), 
        .GT_TXPHINIT                    (sync_txphinit[i]),   
        .GT_TXDLYBYPASS                 (sync_txdlybypass[i]),  
        .GT_TXDLYSRESET                 (sync_txdlysreset[i]),
        .GT_TXDLYEN                     (sync_txdlyen[i]),      
                                     
        .GT_TXDLYSRESETDONE             (gt_txdlysresetdone[i]),
        .GT_TXPHINITDONE                (gt_txphinitdone[i]),  
        .GT_TXPHALIGNDONE               (gt_txphaligndone[i]), 
        
        .GT_TXPHDLYRESET                (sync_txphdlyreset[i]),
        .GT_TXSYNCMODE                  (i == 0),           // GTH, GTP
        .GT_TXSYNCIN                    (gt_txsyncout[0]),  // GTH, GTP
        .GT_TXSYNCALLIN                 (txsyncallin),      // GTH, GTP
        
        .GT_TXSYNCOUT                   (gt_txsyncout[i]),  // GTH, GTP
        .GT_TXSYNCDONE                  (gt_txsyncdone[i]), // GTH, GTP
        
        //---------- GT RX Sync Ports ----------------------
        .GT_RXPHALIGN                   (sync_rxphalign[i]),
        .GT_RXPHALIGNEN                 (sync_rxphalignen[i]),  
        .GT_RXDLYBYPASS                 (sync_rxdlybypass[i]),         
        .GT_RXDLYSRESET                 (sync_rxdlysreset[i]),
        .GT_RXDLYEN                     (sync_rxdlyen[i]),
        .GT_RXDDIEN                     (sync_rxddien[i]),
                                     
        .GT_RXDLYSRESETDONE             (gt_rxdlysresetdone[i]),
        .GT_RXPHALIGNDONE               (gt_rxphaligndone[i]),
                                                                   
        .GT_RXSYNCMODE                  (i == 0),           // GTH                                                                      
        .GT_RXSYNCIN                    (gt_rxsyncout[0]),  // GTH                                                                      
        .GT_RXSYNCALLIN                 (rxsyncallin),      // GTH     
                    
        .GT_RXSYNCOUT                   (gt_rxsyncout[i]),  // GTH  
        .GT_RXSYNCDONE                  (gt_rxsyncdone[i]), // GTH      
                                                                         
        //---------- GT Comma Alignment Ports --------------
        .GT_RXSLIDE                     (PIPE_RXSLIDE[i]),
    
        .GT_RXCOMMADET                  (gt_rxcommadet[i]),                        
        .GT_RXCHARISCOMMA               (gt_rxchariscomma[(4*i)+3:(4*i)]),                      
        .GT_RXBYTEISALIGNED             (gt_rxbyteisaligned[i]),                   
        .GT_RXBYTEREALIGN               (gt_rxbyterealign[i]),
    
        //---------- GT Channel Bonding Ports --------------
        .GT_RXCHANISALIGNED             (PIPE_RXCHANISALIGNED[i]),
        .GT_RXCHBONDEN                  (rxchbonden[i]),
        .GT_RXCHBONDI                   (gt_rxchbondi[i]),
        .GT_RXCHBONDLEVEL               (gt_rxchbondlevel[(3*i)+2:(3*i)]),
        .GT_RXCHBONDMASTER              (rxchbondmaster[i]),
        .GT_RXCHBONDSLAVE               (rxchbondslave[i]),
        .GT_RXCHBONDO                   (gt_rxchbondo[i+1]),
        
        //---------- GT PRBS/Loopback Ports ----------------
        .GT_TXPRBSSEL                   (PIPE_TXPRBSSEL),
        .GT_RXPRBSSEL                   (PIPE_RXPRBSSEL),
        .GT_TXPRBSFORCEERR              (PIPE_TXPRBSFORCEERR),
        .GT_RXPRBSCNTRESET              (PIPE_RXPRBSCNTRESET),
        .GT_LOOPBACK                    (PIPE_LOOPBACK),    
        
        .GT_RXPRBSERR                   (PIPE_RXPRBSERR[i]),
        
        //---------- GT Debug Port -------------------------
        .GT_DMONITOROUT                 (PIPE_DMONITOROUT[(15*i)+14:(15*i)])
    );
    

    
    //---------- GT Wrapper Assignments ----------------------------------------     
    assign oobclk[i]         = (PCIE_OOBCLK_MODE == 1) ? user_oobclk[i] : clk_oobclk;
    
    //---------- Channel Bonding Master Slave Enable ---------------------------
    if (PCIE_CHAN_BOND_EN == "FALSE") 
        begin : channel_bonding_ms_disable
        assign rxchbonden[i]     = 1'd0; 
        assign rxchbondmaster[i] = 1'd0;
        assign rxchbondslave[i]  = 1'd0;
        end 
    else 
        begin : channel_bonding_ms_enable
        assign rxchbonden[i]     = (PCIE_LANE > 1) && (PCIE_CHAN_BOND_EN == "TRUE") ? !rate_gen3[i] : 1'd0; 
        assign rxchbondmaster[i] =  rate_gen3[i] ? 1'd0 : (i == 0);
        assign rxchbondslave[i]  =  rate_gen3[i] ? 1'd0 : (i  > 0);
        end
    
    //---------- Channel Bonding Input Connection ------------------------------
    if (PCIE_CHAN_BOND_EN == "FALSE") 
        begin : channel_bonding_in_disable
        assign gt_rxchbondi[i]                 = 5'd0; 
        assign gt_rxchbondlevel[(3*i)+2:(3*i)] = 3'd0;
        end
    else
        begin : channel_bonding_in_enable
        
        //---------- Channel Bonding (2: Binary-Tree) --------------------------
        if (PCIE_CHAN_BOND == 2) 
        
            begin : channel_bonding_a
            
            case (i)
            
            //---------- Lane 0 --------------------------------
            0 : 
                begin
                assign gt_rxchbondi[0]         = gt_rxchbondo[0];
                assign gt_rxchbondlevel[2:0]   = (PCIE_LANE == 4'd8) ? 3'd4 : 
                                                 (PCIE_LANE >  4'd5) ? 3'd3 : 
                                                 (PCIE_LANE >  4'd3) ? 3'd2 : 
                                                 (PCIE_LANE >  4'd1) ? 3'd1 : 3'd0; 
                end
            //---------- Lane 1 --------------------------------    
            1 : 
                begin
                assign gt_rxchbondi[1]         = gt_rxchbondo[1];
                assign gt_rxchbondlevel[5:3]   = (PCIE_LANE == 4'd8) ? 3'd3 : 
                                                 (PCIE_LANE >  4'd5) ? 3'd2 : 
                                                 (PCIE_LANE >  4'd3) ? 3'd1 : 3'd0; 
                end
            //---------- Lane 2 --------------------------------
            2 : 
                begin
                assign gt_rxchbondi[2]         = gt_rxchbondo[1];
                assign gt_rxchbondlevel[8:6]   = (PCIE_LANE == 4'd8) ? 3'd3 : 
                                                 (PCIE_LANE >  4'd5) ? 3'd2 : 
                                                 (PCIE_LANE >  4'd3) ? 3'd1 : 3'd0; 
                end
            //---------- Lane 3 --------------------------------
            3 : 
                begin
                assign gt_rxchbondi[3]         = gt_rxchbondo[3];
                assign gt_rxchbondlevel[11:9]  = (PCIE_LANE == 4'd8) ? 3'd2 : 
                                                 (PCIE_LANE >  4'd5) ? 3'd1 : 3'd0;
                end
            //---------- Lane 4 --------------------------------
            4 : 
                begin
                assign gt_rxchbondi[4]         = gt_rxchbondo[3];
                assign gt_rxchbondlevel[14:12] = (PCIE_LANE == 4'd8) ? 3'd2 : 
                                                 (PCIE_LANE >  4'd5) ? 3'd1 : 3'd0;
                end
            //---------- Lane 5 --------------------------------
            5 : 
                begin
                assign gt_rxchbondi[5]         = gt_rxchbondo[5];
                assign gt_rxchbondlevel[17:15] = (PCIE_LANE == 4'd8) ? 3'd1 : 3'd0;
                end
            //---------- Lane 6 --------------------------------
            6 : 
                begin
                assign gt_rxchbondi[6]         = gt_rxchbondo[5];
                assign gt_rxchbondlevel[20:18] = (PCIE_LANE == 4'd8) ? 3'd1 : 3'd0;
                end
            //---------- Lane 7 --------------------------------
            7 : 
                begin
                assign gt_rxchbondi[7]         = gt_rxchbondo[7]; 
                assign gt_rxchbondlevel[23:21] = 3'd0;
                end     
            //---------- Default -------------------------------
            default :
                begin
                assign gt_rxchbondi[i]                 = gt_rxchbondo[7]; 
                assign gt_rxchbondlevel[(3*i)+2:(3*i)] = 3'd0;
                end
                
            endcase    
                
            end
            
        //---------- Channel Bonding (0: One-Hop, 1: Daisy Chain) --------------    
        else 
        
            begin : channel_bonding_b
            assign gt_rxchbondi[i]                 = (PCIE_CHAN_BOND == 1) ? gt_rxchbondo[i] : ((i == 0) ? gt_rxchbondo[0] : gt_rxchbondo[1]);
            assign gt_rxchbondlevel[(3*i)+2:(3*i)] = (PCIE_CHAN_BOND == 1) ? (PCIE_LANE-1)-i  : ((PCIE_LANE > 1) && (i == 0));       
            end
        
        end 
        
        end

endgenerate 



//---------- PIPE Wrapper Output -----------------------------------------------
assign PIPE_TXEQ_FS      = 0;//TXEQ_FS;
assign PIPE_TXEQ_LF      = 0;//TXEQ_LF;
assign PIPE_RXELECIDLE   = gt_rxelecidle;
assign PIPE_RXSTATUS     = gt_rxstatus;

assign PIPE_RXDISPERR       = gt_rxdisperr;  
assign PIPE_RXNOTINTABLE    = gt_rxnotintable;
assign PIPE_RXPMARESETDONE  = gt_rxpmaresetdone;
assign PIPE_RXBUFSTATUS     = gt_rxbufstatus;
assign PIPE_TXPHALIGNDONE   = gt_txphaligndone;
assign PIPE_TXPHINITDONE    = gt_txphinitdone;
assign PIPE_TXDLYSRESETDONE = gt_txdlysresetdone;
assign PIPE_RXPHALIGNDONE   = gt_rxphaligndone;
assign PIPE_RXDLYSRESETDONE = gt_rxdlysresetdone;
assign PIPE_RXSYNCDONE      = gt_rxsyncdone;
assign PIPE_RXCOMMADET      = gt_rxcommadet;
assign PIPE_QPLL_LOCK       = qpll_qplllock;
assign PIPE_CPLL_LOCK       = gt_cplllock;   

assign PIPE_PCLK         = clk_pclk;
assign PIPE_PCLK_LOCK    = clk_mmcm_lock; 
assign PIPE_RXCDRLOCK    = 0;//user_rxcdrlock;
assign PIPE_RXUSRCLK     = 0;//clk_rxusrclk; 
assign PIPE_RXOUTCLK     = 0;//clk_rxoutclk;
assign PIPE_TXSYNC_DONE  = 0;//sync_txsync_done;
assign PIPE_RXSYNC_DONE  = 0;//sync_rxsync_done;
assign PIPE_ACTIVE_LANE  = 0;//user_active_lane;
             
assign PIPE_TXOUTCLK_OUT = gt_txoutclk[0];
assign PIPE_RXOUTCLK_OUT = gt_rxoutclk;
assign PIPE_PCLK_SEL_OUT = rate_pclk_sel;
assign PIPE_GEN3_OUT     = rate_gen3[0];

assign PIPE_RXEQ_CONVERGE   = user_rx_converge;
assign PIPE_RXEQ_ADAPT_DONE = (PCIE_GT_DEVICE == "GTP") ? {PCIE_LANE{1'd0}} : eq_rxeq_adapt_done;

assign PIPE_EYESCANDATAERROR = gt_eyescandataerror;
assign PIPE_RST_FSM      = rst_fsm;
assign PIPE_QRST_FSM     = qrst_fsm;
assign PIPE_RATE_FSM     = rate_fsm;
assign PIPE_SYNC_FSM_TX  = sync_fsm_tx;
assign PIPE_SYNC_FSM_RX  = sync_fsm_rx;
assign PIPE_DRP_FSM      = drp_fsm;   
assign PIPE_QDRP_FSM     = 0;//qdrp_fsm;
                        
assign PIPE_RST_IDLE     = &rst_idle;
assign PIPE_QRST_IDLE    = &qrst_idle;
assign PIPE_RATE_IDLE    = &rate_idle;

assign EXT_CH_GT_DRPDO   =  gt_do[(PCIE_LANE*16)-1:0];
assign EXT_CH_GT_DRPRDY  =  gt_rdy[(PCIE_LANE-1):0];
assign EXT_CH_GT_DRPCLK  =  clk_dclk;

assign PIPE_DEBUG_0      = (PCIE_DEBUG_MODE == 1) ? gt_txresetdone                  : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_1      = (PCIE_DEBUG_MODE == 1) ? gt_rxresetdone                  : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_2      = (PCIE_DEBUG_MODE == 1) ? gt_phystatus                    : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_3      = (PCIE_DEBUG_MODE == 1) ? gt_rxvalid                      : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_4      = (PCIE_DEBUG_MODE == 1) ? clk_dclk                        : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_5      = (PCIE_DEBUG_MODE == 1) ? drp_mux_en                      : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_6      = (PCIE_DEBUG_MODE == 1) ? drp_mux_we                      : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_7      = (PCIE_DEBUG_MODE == 1) ? gt_rdy                          : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_8      = (PCIE_DEBUG_MODE == 1) ? user_rx_converge                : {PCIE_LANE{1'b0}};
assign PIPE_DEBUG_9      = (PCIE_DEBUG_MODE == 1) ? PIPE_TXELECIDLE                 : {PCIE_LANE{1'b0}};

assign PIPE_DEBUG[ 1:0]  = (PCIE_DEBUG_MODE == 1) ? PIPE_TXEQ_CONTROL[1:0] : 2'd0;
assign PIPE_DEBUG[ 5:2]  = (PCIE_DEBUG_MODE == 1) ? PIPE_TXEQ_PRESET[3:0]  : 4'd0;
assign PIPE_DEBUG[31:6]  = 26'd0;



endmodule


`timescale 1ns/1ps
module model_ap2_tst_gtp_pipe_reset #
(

    //---------- Global ------------------------------------
    parameter PCIE_SIM_SPEEDUP = "FALSE",                   // PCIe sim speedup 
    parameter PCIE_LANE        = 1,                         // PCIe number of lanes
    //---------- Local -------------------------------------
    parameter CFG_WAIT_MAX     = 6'd63,                     // Configuration wait max
    parameter BYPASS_RXCDRLOCK = 1                          // Bypass RXCDRLOCK

)

(

    //---------- Input -------------------------------------
    input                           RST_CLK,
    input                           RST_RXUSRCLK,
    input                           RST_DCLK,
    input                           RST_RST_N,
    input       [PCIE_LANE-1:0]     RST_DRP_DONE,
    input       [PCIE_LANE-1:0]     RST_RXPMARESETDONE,
    input                           RST_PLLLOCK,
    input       [PCIE_LANE-1:0]     RST_RATE_IDLE,
    input       [PCIE_LANE-1:0]     RST_RXCDRLOCK,
    input                           RST_MMCM_LOCK,
    input       [PCIE_LANE-1:0]     RST_RESETDONE,
    input       [PCIE_LANE-1:0]     RST_PHYSTATUS,
    input       [PCIE_LANE-1:0]     RST_TXSYNC_DONE,
    
    //---------- Output ------------------------------------
    output                          RST_CPLLRESET,
    output                          RST_CPLLPD,
    output reg                      RST_DRP_START,
    output reg                      RST_DRP_X16,
    output                          RST_RXUSRCLK_RESET,
    output                          RST_DCLK_RESET,
    output                          RST_GTRESET,
    output                          RST_USERRDY,
    output                          RST_TXSYNC_START,
    output                          RST_IDLE,
    output      [ 4:0]              RST_FSM

);

    //---------- Input Register ----------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     drp_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxpmaresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             plllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rate_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxcdrlock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     resetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     phystatus_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     txsync_done_reg1;  
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     drp_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxpmaresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             plllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rate_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxcdrlock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     resetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     phystatus_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     txsync_done_reg2;
    
    //---------- Internal Signal ---------------------------
    reg         [ 5:0]              cfg_wait_cnt      =  6'd0;
    
    //---------- Output Register ---------------------------
    reg                             pllreset          =  1'd0;
    reg                             pllpd             =  1'd0;
    reg                             rxusrclk_rst_reg1 =  1'd0;
    reg                             rxusrclk_rst_reg2 =  1'd0;
    reg                             dclk_rst_reg1     =  1'd0;
    reg                             dclk_rst_reg2     =  1'd0;
    reg                             gtreset           =  1'd0;
    reg                             userrdy           =  1'd0;
    reg         [ 4:0]              fsm               =  5'h1;                 
   
    //---------- FSM ---------------------------------------                                         
    localparam                      FSM_IDLE             = 5'h0; 
    localparam                      FSM_CFG_WAIT         = 5'h1;
    localparam                      FSM_PLLRESET         = 5'h2; 
    localparam                      FSM_DRP_X16_START    = 5'h3;
    localparam                      FSM_DRP_X16_DONE     = 5'h4;   
    localparam                      FSM_PLLLOCK          = 5'h5;
    localparam                      FSM_GTRESET          = 5'h6;
    localparam                      FSM_RXPMARESETDONE_1 = 5'h7; 
    localparam                      FSM_RXPMARESETDONE_2 = 5'h8; 
    localparam                      FSM_DRP_X20_START    = 5'h9;
    localparam                      FSM_DRP_X20_DONE     = 5'hA;                    
    localparam                      FSM_MMCM_LOCK        = 5'hB;  
    localparam                      FSM_RESETDONE        = 5'hC;  
    localparam                      FSM_TXSYNC_START     = 5'hD;
    localparam                      FSM_TXSYNC_DONE      = 5'hE;                                 

    

//---------- Input FF ----------------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------  
        drp_done_reg1       <= {PCIE_LANE{1'd0}};   
        rxpmaresetdone_reg1 <= {PCIE_LANE{1'd0}}; 
        plllock_reg1        <= 1'd0; 
        rate_idle_reg1      <= {PCIE_LANE{1'd0}}; 
        rxcdrlock_reg1      <= {PCIE_LANE{1'd0}}; 
        mmcm_lock_reg1      <= 1'd0; 
        resetdone_reg1      <= {PCIE_LANE{1'd0}}; 
        phystatus_reg1      <= {PCIE_LANE{1'd0}}; 
        txsync_done_reg1    <= {PCIE_LANE{1'd0}}; 
        //---------- 2nd Stage FF --------------------------
        drp_done_reg2       <= {PCIE_LANE{1'd0}};
        rxpmaresetdone_reg2 <= {PCIE_LANE{1'd0}}; 
        plllock_reg2        <= 1'd0; 
        rate_idle_reg2      <= {PCIE_LANE{1'd0}}; 
        rxcdrlock_reg2      <= {PCIE_LANE{1'd0}}; 
        mmcm_lock_reg2      <= 1'd0;
        resetdone_reg2      <= {PCIE_LANE{1'd0}}; 
        phystatus_reg2      <= {PCIE_LANE{1'd0}}; 
        txsync_done_reg2    <= {PCIE_LANE{1'd0}}; 
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------   
        drp_done_reg1       <= RST_DRP_DONE; 
        rxpmaresetdone_reg1 <= RST_RXPMARESETDONE; 
        plllock_reg1        <= RST_PLLLOCK;
        rate_idle_reg1      <= RST_RATE_IDLE;
        rxcdrlock_reg1      <= RST_RXCDRLOCK;
        mmcm_lock_reg1      <= RST_MMCM_LOCK;
        resetdone_reg1      <= RST_RESETDONE;
        phystatus_reg1      <= RST_PHYSTATUS;
        txsync_done_reg1    <= RST_TXSYNC_DONE;
        //---------- 2nd Stage FF --------------------------
        drp_done_reg2       <= drp_done_reg1;
        rxpmaresetdone_reg2 <= rxpmaresetdone_reg1;
        plllock_reg2        <= plllock_reg1;
        rate_idle_reg2      <= rate_idle_reg1;
        rxcdrlock_reg2      <= rxcdrlock_reg1;
        mmcm_lock_reg2      <= mmcm_lock_reg1;
        resetdone_reg2      <= resetdone_reg1;
        phystatus_reg2      <= phystatus_reg1;
        txsync_done_reg2    <= txsync_done_reg1;   
        end
        
end    



//---------- Configuration Reset Wait Counter ----------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        cfg_wait_cnt <= 6'd0;
    else
    
        //---------- Increment Configuration Reset Wait Counter
        if ((fsm == FSM_CFG_WAIT) && (cfg_wait_cnt < CFG_WAIT_MAX))
            cfg_wait_cnt <= cfg_wait_cnt + 6'd1;
            
        //---------- Hold Configuration Reset Wait Counter -
        else if ((fsm == FSM_CFG_WAIT) && (cfg_wait_cnt == CFG_WAIT_MAX))
            cfg_wait_cnt <= cfg_wait_cnt;
            
        //---------- Reset Configuration Reset Wait Counter 
        else
            cfg_wait_cnt <= 6'd0;
        
end 



//---------- PIPE Reset FSM ----------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        begin
        fsm      <= FSM_CFG_WAIT;
        pllreset <= 1'd0;
        pllpd    <= 1'd0;
        gtreset  <= 1'd0;
        userrdy  <= 1'd0;
        end
    else
        begin
        
        case (fsm)
            
        //---------- Idle State ----------------------------
        FSM_IDLE :
        
            begin
            if (!RST_RST_N)
                begin
                fsm      <= FSM_CFG_WAIT;
                pllreset <= 1'd0;
                pllpd    <= 1'd0;
                gtreset  <= 1'd0;
                userrdy  <= 1'd0;
                end
            else
                begin
                fsm      <= FSM_IDLE;
                pllreset <= pllreset;
                pllpd    <= pllpd;
                gtreset  <= gtreset;
                userrdy  <= userrdy;
                end
            end  
            
        //----------  Wait for Configuration Reset Delay ---
        FSM_CFG_WAIT :
          
            begin
            fsm       <= ((cfg_wait_cnt == CFG_WAIT_MAX) ? FSM_PLLRESET : FSM_CFG_WAIT);
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end 
            
        //---------- Hold PLL and GTP Channel in Reset ----
        FSM_PLLRESET :
        
            begin
            fsm       <= (((~plllock_reg2) && (&(~resetdone_reg2))) ? FSM_DRP_X16_START : FSM_PLLRESET);
            pllreset  <= 1'd1;
            pllpd     <= pllpd;
            gtreset   <= 1'd1;
            userrdy   <= userrdy;
            end  

        //---------- Start DRP x16 -------------------------
        FSM_DRP_X16_START :
            
            begin
            fsm       <= &(~drp_done_reg2) ? FSM_DRP_X16_DONE : FSM_DRP_X16_START;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for DRP x16 Done -----------------    
        FSM_DRP_X16_DONE :
        
            begin  
            fsm       <= (&drp_done_reg2) ? FSM_PLLLOCK : FSM_DRP_X16_DONE;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  

        //---------- Wait for PLL Lock --------------------
        FSM_PLLLOCK :
        
            begin
            fsm       <= (plllock_reg2 ? FSM_GTRESET : FSM_PLLLOCK);
            pllreset  <= 1'd0;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end

        //---------- Release GTRESET -----------------------
        FSM_GTRESET :
        
            begin
            fsm       <= FSM_RXPMARESETDONE_1;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= 1'b0;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for RXPMARESETDONE Assertion -----  
        FSM_RXPMARESETDONE_1 :
        
            begin
            fsm       <= (&rxpmaresetdone_reg2 || (PCIE_SIM_SPEEDUP == "TRUE")) ? FSM_RXPMARESETDONE_2 : FSM_RXPMARESETDONE_1;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  

        //---------- Wait for RXPMARESETDONE De-assertion --
        FSM_RXPMARESETDONE_2 :
        
            begin
            fsm       <= (&(~rxpmaresetdone_reg2) || (PCIE_SIM_SPEEDUP == "TRUE")) ? FSM_DRP_X20_START : FSM_RXPMARESETDONE_2;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  
            
        //---------- Start DRP x20 -------------------------
        FSM_DRP_X20_START :
            
            begin
            fsm       <= &(~drp_done_reg2) ? FSM_DRP_X20_DONE : FSM_DRP_X20_START;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for DRP x20 Done -----------------    
        FSM_DRP_X20_DONE :
        
            begin  
            fsm       <= (&drp_done_reg2) ? FSM_MMCM_LOCK : FSM_DRP_X20_DONE;
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end      

        //---------- Wait for MMCM and RX CDR Lock ---------
        FSM_MMCM_LOCK :
        
            begin  
            if (mmcm_lock_reg2 && (&rxcdrlock_reg2 || (BYPASS_RXCDRLOCK == 1)))
                begin
                fsm       <= FSM_RESETDONE;
                pllreset  <= pllreset;
                pllpd     <= pllpd;
                gtreset   <= gtreset;
                userrdy   <= 1'd1;
                end
            else
                begin
                fsm       <= FSM_MMCM_LOCK;
                pllreset  <= pllreset;
                pllpd     <= pllpd;
                gtreset   <= gtreset;
                userrdy   <= 1'd0;
                end
            end

        //---------- Wait for [TX/RX]RESETDONE and PHYSTATUS 
        FSM_RESETDONE :
        
            begin
            fsm       <= (&resetdone_reg2 && (&(~phystatus_reg2)) ? FSM_TXSYNC_START : FSM_RESETDONE);  
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Start TX Sync -------------------------
        FSM_TXSYNC_START :
        
            begin
            fsm       <= (&(~txsync_done_reg2) ? FSM_TXSYNC_DONE : FSM_TXSYNC_START);
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for TX Sync Done -----------------
        FSM_TXSYNC_DONE :
        
            begin
            fsm       <= (&txsync_done_reg2 ? FSM_IDLE : FSM_TXSYNC_DONE);
            pllreset  <= pllreset;
            pllpd     <= pllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end     
            
        //---------- Default State -------------------------
        default :
        
            begin
            fsm       <= FSM_CFG_WAIT;
            pllreset  <= 1'd0;
            pllpd     <= 1'd0;
            gtreset   <= 1'd0;
            userrdy   <= 1'd0;
            end

        endcase
        
        end
        
end



//---------- RXUSRCLK Reset Synchronizer ---------------------------------------
always @ (posedge RST_RXUSRCLK)
begin

    if (pllreset) 
        begin
        rxusrclk_rst_reg1 <= 1'd1;
        rxusrclk_rst_reg2 <= 1'd1;
        end
    else
        begin
        rxusrclk_rst_reg1 <= 1'd0;
        rxusrclk_rst_reg2 <= rxusrclk_rst_reg1;
        end   
          
end  

//---------- DCLK Reset Synchronizer -------------------------------------------
always @ (posedge RST_DCLK)
begin

    if (fsm == FSM_CFG_WAIT)
        begin
        dclk_rst_reg1 <= 1'd1;
        dclk_rst_reg2 <= dclk_rst_reg1;
        end
    else
        begin
        dclk_rst_reg1 <= 1'd0;
        dclk_rst_reg2 <= dclk_rst_reg1;
        end   
          
end  



//---------- PIPE Reset Output -------------------------------------------------
assign RST_CPLLRESET      = pllreset;
assign RST_CPLLPD         = pllpd;
assign RST_RXUSRCLK_RESET = rxusrclk_rst_reg2;
assign RST_DCLK_RESET     = dclk_rst_reg2;
assign RST_GTRESET        = gtreset;  
assign RST_USERRDY        = userrdy;
assign RST_TXSYNC_START   = (fsm == FSM_TXSYNC_START);
assign RST_IDLE           = (fsm == FSM_IDLE);
assign RST_FSM            = fsm;                   



//--------------------------------------------------------------------------------------------------
//  Register Output
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N) 
        begin
        RST_DRP_START <= 1'd0;
        RST_DRP_X16   <= 1'd0;
        end
    else
        begin
        RST_DRP_START <= (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X20_START); 
        RST_DRP_X16   <= (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X16_DONE);
        end
        
end  



endmodule


`timescale 1ns/1ps
module model_ap2_tst_pipe_reset #
(

    //---------- Global ------------------------------------
    parameter PCIE_SIM_SPEEDUP  = "FALSE",                  // PCIe sim speedup
    parameter PCIE_GT_DEVICE    = "GTX",
    parameter PCIE_PLL_SEL      = "CPLL",                   // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_POWER_SAVING = "TRUE",                   // PCIe power saving
    parameter PCIE_TXBUF_EN     = "FALSE",                  // PCIe TX buffer enable
    parameter PCIE_LANE         = 1,                        // PCIe number of lanes
    //---------- Local -------------------------------------
    parameter CFG_WAIT_MAX      = 6'd63,                    // Configuration wait max
    parameter BYPASS_RXCDRLOCK  = 1                         // Bypass RXCDRLOCK

)

(

    //---------- Input -------------------------------------
    input                           RST_CLK,
    input                           RST_RXUSRCLK,
    input                           RST_DCLK,
    input                           RST_RST_N,
    input       [PCIE_LANE-1:0]     RST_DRP_DONE,
    input       [PCIE_LANE-1:0]     RST_RXPMARESETDONE,
    input       [PCIE_LANE-1:0]     RST_CPLLLOCK,
    input                           RST_QPLL_IDLE,
    input       [PCIE_LANE-1:0]     RST_RATE_IDLE,
    input       [PCIE_LANE-1:0]     RST_RXCDRLOCK,
    input                           RST_MMCM_LOCK,
    input       [PCIE_LANE-1:0]     RST_RESETDONE,
    input       [PCIE_LANE-1:0]     RST_PHYSTATUS,
    input       [PCIE_LANE-1:0]     RST_TXSYNC_DONE,
    
    //---------- Output ------------------------------------
    output                          RST_CPLLRESET,
    output                          RST_CPLLPD,
    output reg                      RST_DRP_START,
    output reg                      RST_DRP_X16X20_MODE,
    output reg                      RST_DRP_X16,
    output                          RST_RXUSRCLK_RESET,
    output                          RST_DCLK_RESET,
    output                          RST_GTRESET,
    output                          RST_USERRDY,
    output                          RST_TXSYNC_START,
    output                          RST_IDLE,
    output      [4:0]               RST_FSM

);

    //---------- Input Register ----------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     drp_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxpmaresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     cplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             qpll_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rate_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxcdrlock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     resetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     phystatus_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     txsync_done_reg1;  
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     drp_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxpmaresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     cplllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             qpll_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rate_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     rxcdrlock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     resetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     phystatus_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     txsync_done_reg2;
    
    //---------- Internal Signal ---------------------------
    reg         [ 5:0]              cfg_wait_cnt      =  6'd0;
    
    //---------- Output Register ---------------------------
    reg                             cpllreset         =  1'd0;
    reg                             cpllpd            =  1'd0;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             rxusrclk_rst_reg1 =  1'd0;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             rxusrclk_rst_reg2 =  1'd0;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             dclk_rst_reg1     =  1'd0;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             dclk_rst_reg2     =  1'd0;
    reg                             gtreset           =  1'd0;
    reg                             userrdy           =  1'd0;
    reg         [4:0]               fsm               =  5'h2;
   
    //---------- FSM ---------------------------------------                                         
    localparam                      FSM_IDLE             = 5'h0;
    localparam                      FSM_CFG_WAIT         = 5'h1;
    localparam                      FSM_CPLLRESET        = 5'h2;
    localparam                      FSM_DRP_X16_START    = 5'h3;
    localparam                      FSM_DRP_X16_DONE     = 5'h4;
    localparam                      FSM_CPLLLOCK         = 5'h5;
    localparam                      FSM_DRP              = 5'h6;
    localparam                      FSM_GTRESET          = 5'h7;
    localparam                      FSM_RXPMARESETDONE_1 = 5'h8;
    localparam                      FSM_RXPMARESETDONE_2 = 5'h9;
    localparam                      FSM_DRP_X20_START    = 5'hA;
    localparam                      FSM_DRP_X20_DONE     = 5'hB;
    localparam                      FSM_MMCM_LOCK        = 5'hC;
    localparam                      FSM_RESETDONE        = 5'hD;
    localparam                      FSM_CPLL_PD          = 5'hE;
    localparam                      FSM_TXSYNC_START     = 5'hF;
    localparam                      FSM_TXSYNC_DONE      = 5'h10;

    

//---------- Input FF ----------------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------    
        drp_done_reg1       <= {PCIE_LANE{1'd0}};   
        rxpmaresetdone_reg1 <= {PCIE_LANE{1'd0}}; 
        cplllock_reg1       <= {PCIE_LANE{1'd0}}; 
        qpll_idle_reg1      <= 1'd0;
        rate_idle_reg1      <= {PCIE_LANE{1'd0}}; 
        rxcdrlock_reg1      <= {PCIE_LANE{1'd0}}; 
        mmcm_lock_reg1      <= 1'd0; 
        resetdone_reg1      <= {PCIE_LANE{1'd0}}; 
        phystatus_reg1      <= {PCIE_LANE{1'd0}}; 
        txsync_done_reg1    <= {PCIE_LANE{1'd0}}; 
        //---------- 2nd Stage FF --------------------------
        drp_done_reg2       <= {PCIE_LANE{1'd0}};
        rxpmaresetdone_reg2 <= {PCIE_LANE{1'd0}}; 
        cplllock_reg2       <= {PCIE_LANE{1'd0}}; 
        qpll_idle_reg2      <= 1'd0;
        rate_idle_reg2      <= {PCIE_LANE{1'd0}}; 
        rxcdrlock_reg2      <= {PCIE_LANE{1'd0}}; 
        mmcm_lock_reg2      <= 1'd0;
        resetdone_reg2      <= {PCIE_LANE{1'd0}}; 
        phystatus_reg2      <= {PCIE_LANE{1'd0}}; 
        txsync_done_reg2    <= {PCIE_LANE{1'd0}}; 
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------  
        drp_done_reg1       <= RST_DRP_DONE; 
        rxpmaresetdone_reg1 <= RST_RXPMARESETDONE;   
        cplllock_reg1       <= RST_CPLLLOCK;
        qpll_idle_reg1      <= RST_QPLL_IDLE;
        rate_idle_reg1      <= RST_RATE_IDLE;
        rxcdrlock_reg1      <= RST_RXCDRLOCK;
        mmcm_lock_reg1      <= RST_MMCM_LOCK;
        resetdone_reg1      <= RST_RESETDONE;
        phystatus_reg1      <= RST_PHYSTATUS;
        txsync_done_reg1    <= RST_TXSYNC_DONE;
        //---------- 2nd Stage FF --------------------------
        drp_done_reg2       <= drp_done_reg1;
        rxpmaresetdone_reg2 <= rxpmaresetdone_reg1;
        cplllock_reg2       <= cplllock_reg1;
        qpll_idle_reg2      <= qpll_idle_reg1;
        rate_idle_reg2      <= rate_idle_reg1;
        rxcdrlock_reg2      <= rxcdrlock_reg1;
        mmcm_lock_reg2      <= mmcm_lock_reg1;
        resetdone_reg2      <= resetdone_reg1;
        phystatus_reg2      <= phystatus_reg1;
        txsync_done_reg2    <= txsync_done_reg1;   
        end
        
end    



//---------- Configuration Reset Wait Counter ----------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        cfg_wait_cnt <= 6'd0;
    else
    
        //---------- Increment Configuration Reset Wait Counter
        if ((fsm == FSM_CFG_WAIT) && (cfg_wait_cnt < CFG_WAIT_MAX))
            cfg_wait_cnt <= cfg_wait_cnt + 6'd1;
            
        //---------- Hold Configuration Reset Wait Counter -
        else if ((fsm == FSM_CFG_WAIT) && (cfg_wait_cnt == CFG_WAIT_MAX))
            cfg_wait_cnt <= cfg_wait_cnt;
            
        //---------- Reset Configuration Reset Wait Counter 
        else
            cfg_wait_cnt <= 6'd0;
        
end 



//---------- PIPE Reset FSM ----------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N)
        begin
        fsm       <= FSM_CFG_WAIT;
        cpllreset <= 1'd0;
        cpllpd    <= 1'd0;
        gtreset   <= 1'd0;
        userrdy   <= 1'd0;
        end
    else
        begin
        
        case (fsm)
            
        //---------- Idle State ----------------------------
        FSM_IDLE :
        
            begin
            if (!RST_RST_N)
                begin
                fsm       <= FSM_CFG_WAIT;
                cpllreset <= 1'd0;
                cpllpd    <= 1'd0;
                gtreset   <= 1'd0;
                userrdy   <= 1'd0;
                end
            else
                begin
                fsm       <= FSM_IDLE;
                cpllreset <= cpllreset;
                cpllpd    <= cpllpd;
                gtreset   <= gtreset;
                userrdy   <= userrdy;
                end
            end  
            
        //----------  Wait for Configuration Reset Delay ---
        FSM_CFG_WAIT :
          
            begin
            fsm       <= ((cfg_wait_cnt == CFG_WAIT_MAX) ? FSM_CPLLRESET : FSM_CFG_WAIT);
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end 
            
        //---------- Hold CPLL and GTX Channel in Reset ----
        FSM_CPLLRESET :
        
            begin
            fsm       <= ((&(~cplllock_reg2) && (&(~resetdone_reg2))) ?  FSM_CPLLLOCK : FSM_CPLLRESET);
            cpllreset <= 1'd1;
            cpllpd    <= cpllpd;
            gtreset   <= 1'd1;
            userrdy   <= userrdy;
            end  

        //---------- Wait for CPLL Lock --------------------
        FSM_CPLLLOCK :
        
            begin
            fsm       <= (&cplllock_reg2 ? FSM_DRP : FSM_CPLLLOCK);
            cpllreset <= 1'd0;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end

        //---------- Wait for DRP Done to Setup Gen1 -------
        FSM_DRP :
        
            begin
            fsm       <= (&rate_idle_reg2 ? ((PCIE_GT_DEVICE == "GTX") ? FSM_GTRESET : FSM_DRP_X16_START) : FSM_DRP);
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end

        //---------- Start DRP x16 -------------------------
        FSM_DRP_X16_START :
            
            begin
            fsm       <= &(~drp_done_reg2) ? FSM_DRP_X16_DONE : FSM_DRP_X16_START;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for DRP x16 Done -----------------    
        FSM_DRP_X16_DONE :
        
            begin  
            fsm       <= (&drp_done_reg2) ? FSM_GTRESET : FSM_DRP_X16_DONE;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  

        //---------- Release GTX Channel Reset -------------
        FSM_GTRESET :
        
            begin
            fsm       <= (PCIE_GT_DEVICE == "GTX") ? FSM_MMCM_LOCK : FSM_RXPMARESETDONE_1;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= 1'b0;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for RXPMARESETDONE Assertion -----
        FSM_RXPMARESETDONE_1 :
        
            begin
            fsm       <= (&rxpmaresetdone_reg2 || (PCIE_SIM_SPEEDUP == "TRUE")) ? FSM_RXPMARESETDONE_2 : FSM_RXPMARESETDONE_1;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  

        //---------- Wait for RXPMARESETDONE De-assertion --
        FSM_RXPMARESETDONE_2 :
        
            begin
            fsm       <= (&(~rxpmaresetdone_reg2) || (PCIE_SIM_SPEEDUP == "TRUE")) ? FSM_DRP_X20_START : FSM_RXPMARESETDONE_2;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end  
            
        //---------- Start DRP x20 -------------------------
        FSM_DRP_X20_START :
            
            begin
            fsm       <= &(~drp_done_reg2) ? FSM_DRP_X20_DONE : FSM_DRP_X20_START;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for DRP x20 Done -----------------    
        FSM_DRP_X20_DONE :
        
            begin  
            fsm       <= (&drp_done_reg2) ? FSM_MMCM_LOCK : FSM_DRP_X20_DONE;
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end   

        //---------- Wait for MMCM and RX CDR Lock ---------
        FSM_MMCM_LOCK :
        
            begin  
            if (mmcm_lock_reg2 && (&rxcdrlock_reg2 || (BYPASS_RXCDRLOCK == 1)) && (qpll_idle_reg2 || (PCIE_PLL_SEL == "CPLL")))
                begin
                fsm       <= FSM_RESETDONE;
                cpllreset <= cpllreset;
                cpllpd    <= cpllpd;
                gtreset   <= gtreset;
                userrdy   <= 1'd1;
                end
            else
                begin
                fsm       <= FSM_MMCM_LOCK;
                cpllreset <= cpllreset;
                cpllpd    <= cpllpd;
                gtreset   <= gtreset;
                userrdy   <= 1'd0;
                end
            end

        //---------- Wait for [TX/RX]RESETDONE and PHYSTATUS 
        FSM_RESETDONE :
        
            begin
            fsm       <= (&resetdone_reg2 && (&(~phystatus_reg2)) ? FSM_CPLL_PD : FSM_RESETDONE);  
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Power-Down CPLL if QPLL is Used for Gen1/Gen2
        FSM_CPLL_PD :
        
            begin
            fsm       <= ((PCIE_TXBUF_EN == "TRUE") ? FSM_IDLE : FSM_TXSYNC_START);
            cpllreset <= cpllreset;
            cpllpd    <= (PCIE_PLL_SEL == "QPLL");
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
        
        //---------- Start TX Sync -------------------------
        FSM_TXSYNC_START :
        
            begin
            fsm       <= (&(~txsync_done_reg2) ? FSM_TXSYNC_DONE : FSM_TXSYNC_START);
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end
            
        //---------- Wait for TX Sync Done -----------------
        FSM_TXSYNC_DONE :
        
            begin
            fsm       <= (&txsync_done_reg2 ? FSM_IDLE : FSM_TXSYNC_DONE);
            cpllreset <= cpllreset;
            cpllpd    <= cpllpd;
            gtreset   <= gtreset;
            userrdy   <= userrdy;
            end     
            
        //---------- Default State -------------------------
        default :
        
            begin
            fsm       <= FSM_CFG_WAIT;
            cpllreset <= 1'd0;
            cpllpd    <= 1'd0;
            gtreset   <= 1'd0;
            userrdy   <= 1'd0;
            end

        endcase
        
        end
        
end



//---------- RXUSRCLK Reset Synchronizer ---------------------------------------
always @ (posedge RST_RXUSRCLK)
begin

    if (cpllreset) 
        begin
        rxusrclk_rst_reg1 <= 1'd1;
        rxusrclk_rst_reg2 <= 1'd1;
        end
    else
        begin
        rxusrclk_rst_reg1 <= 1'd0;
        rxusrclk_rst_reg2 <= rxusrclk_rst_reg1;
        end   
          
end  



//---------- DCLK Reset Synchronizer -------------------------------------------
always @ (posedge RST_DCLK)
begin

    if (fsm == FSM_CFG_WAIT)
        begin
        dclk_rst_reg1 <= 1'd1;
        dclk_rst_reg2 <= dclk_rst_reg1;
        end
    else
        begin
        dclk_rst_reg1 <= 1'd0;
        dclk_rst_reg2 <= dclk_rst_reg1;
        end   
          
end  



//---------- PIPE Reset Output -------------------------------------------------
assign RST_CPLLRESET       = cpllreset; 
assign RST_CPLLPD          = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : cpllpd);
assign RST_RXUSRCLK_RESET  = rxusrclk_rst_reg2;
assign RST_DCLK_RESET      = dclk_rst_reg2;
assign RST_GTRESET         = gtreset;  
assign RST_USERRDY         = userrdy;
assign RST_TXSYNC_START    = (fsm == FSM_TXSYNC_START);
assign RST_IDLE            = (fsm == FSM_IDLE);
assign RST_FSM             = fsm;                   




//--------------------------------------------------------------------------------------------------
//  Register Output
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_CLK)
begin

    if (!RST_RST_N) 
        begin
        RST_DRP_START       <= 1'd0;
        RST_DRP_X16X20_MODE <= 1'd0; 
        RST_DRP_X16         <= 1'd0;
        end
    else
        begin
        RST_DRP_START       <= (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X20_START); 
        RST_DRP_X16X20_MODE <= (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X16_DONE) || (fsm == FSM_DRP_X20_START) || (fsm == FSM_DRP_X20_DONE);
        RST_DRP_X16         <= (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X16_DONE);
        end
        
end  



endmodule


`timescale 1ns/1ps
module model_ap2_tst_qpll_reset #
(

    //---------- Global ------------------------------------
    parameter PCIE_PLL_SEL       = "CPLL",                  // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_POWER_SAVING  = "TRUE",                  // PCIe power saving
    parameter PCIE_LANE          = 1,                       // PCIe number of lanes
    parameter BYPASS_COARSE_OVRD = 1                        // Bypass coarse frequency override

)

(

    //---------- Input -------------------------------------
    input                           QRST_CLK,
    input                           QRST_RST_N,
    input                           QRST_MMCM_LOCK,
    input       [PCIE_LANE-1:0]     QRST_CPLLLOCK,
    input       [(PCIE_LANE-1)>>2:0]QRST_DRP_DONE,
    input       [(PCIE_LANE-1)>>2:0]QRST_QPLLLOCK,
    input       [ 1:0]              QRST_RATE,
    input       [PCIE_LANE-1:0]     QRST_QPLLRESET_IN,
    input       [PCIE_LANE-1:0]     QRST_QPLLPD_IN,
    
    //---------- Output ------------------------------------                     
    output                          QRST_OVRD,
    output                          QRST_DRP_START,
    output                          QRST_QPLLRESET_OUT,
    output                          QRST_QPLLPD_OUT,
    output                          QRST_IDLE,
    output      [3:0]               QRST_FSM

);

    //---------- Input Register ----------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     cplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [(PCIE_LANE-1)>>2:0]drp_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [(PCIE_LANE-1)>>2:0]qplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]              rate_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     qpllreset_in_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     qpllpd_in_reg1;

(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                             mmcm_lock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     cplllock_reg2;  
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [(PCIE_LANE-1)>>2:0]drp_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [(PCIE_LANE-1)>>2:0]qplllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]              rate_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     qpllreset_in_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0]     qpllpd_in_reg2;
    
    //---------- Output Register  --------------------------
    reg                             ovrd              =  1'd0;
    reg                             qpllreset         =  1'd1;
    reg                             qpllpd            =  1'd0;
    reg         [3:0]               fsm               =  2;                 
   
    //---------- FSM ---------------------------------------                                         
    localparam                      FSM_IDLE          = 1;//12'b000000000001; 
    localparam                      FSM_WAIT_LOCK     = 2;//12'b000000000010;
    localparam                      FSM_MMCM_LOCK     = 3;//12'b000000000100;   
    localparam                      FSM_DRP_START_NOM = 4;//12'b000000001000;
    localparam                      FSM_DRP_DONE_NOM  = 5;//12'b000000010000;
    localparam                      FSM_QPLLLOCK      = 6;//12'b000000100000;
    localparam                      FSM_DRP_START_OPT = 7;//12'b000001000000;                            
    localparam                      FSM_DRP_DONE_OPT  = 8;//12'b000010000000;
    localparam                      FSM_QPLL_RESET    = 9;//12'b000100000000;                                                         
    localparam                      FSM_QPLLLOCK2     = 10;//12'b001000000000;
    localparam                      FSM_QPLL_PDRESET  = 11;//12'b010000000000;
    localparam                      FSM_QPLL_PD       = 12;//12'b100000000000;                                         
 
 
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge QRST_CLK)
begin

    if (!QRST_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------
        mmcm_lock_reg1    <=  1'd0;
        cplllock_reg1     <= {PCIE_LANE{1'd1}}; 
        drp_done_reg1     <= {(((PCIE_LANE-1)>>2)+1){1'd0}};     
        qplllock_reg1     <= {(((PCIE_LANE-1)>>2)+1){1'd0}}; 
        rate_reg1         <=  2'd0; 
        qpllreset_in_reg1 <= {PCIE_LANE{1'd1}}; 
        qpllpd_in_reg1    <= {PCIE_LANE{1'd0}}; 
        //---------- 2nd Stage FF --------------------------
        mmcm_lock_reg2    <=  1'd0;
        cplllock_reg2     <= {PCIE_LANE{1'd1}};
        drp_done_reg2     <= {(((PCIE_LANE-1)>>2)+1){1'd0}}; 
        qplllock_reg2     <= {(((PCIE_LANE-1)>>2)+1){1'd0}}; 
        rate_reg2         <=  2'd0;
        qpllreset_in_reg2 <= {PCIE_LANE{1'd1}}; 
        qpllpd_in_reg2    <= {PCIE_LANE{1'd0}};  
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        mmcm_lock_reg1    <= QRST_MMCM_LOCK;   
        cplllock_reg1     <= QRST_CPLLLOCK; 
        drp_done_reg1     <= QRST_DRP_DONE; 
        qplllock_reg1     <= QRST_QPLLLOCK;
        rate_reg1         <= QRST_RATE; 
        qpllreset_in_reg1 <= QRST_QPLLRESET_IN;
        qpllpd_in_reg1    <= QRST_QPLLPD_IN;
        //---------- 2nd Stage FF --------------------------
        mmcm_lock_reg2    <= mmcm_lock_reg1;
        cplllock_reg2     <= cplllock_reg1;
        drp_done_reg2     <= drp_done_reg1; 
        qplllock_reg2     <= qplllock_reg1;
        rate_reg2         <= rate_reg1;
        qpllreset_in_reg2 <= qpllreset_in_reg1;
        qpllpd_in_reg2    <= qpllpd_in_reg1;
        end
        
end    



//---------- QPLL Reset FSM ----------------------------------------------------
always @ (posedge QRST_CLK)
begin

    if (!QRST_RST_N)
        begin
        fsm       <= FSM_WAIT_LOCK;
        ovrd      <= 1'd0;
        qpllreset <= 1'd1;
        qpllpd    <= 1'd0;
        end
    else
        begin
        
        case (fsm)
            
        //---------- Idle State ----------------------------
        FSM_IDLE :
        
            begin
            if (!QRST_RST_N)
                begin
                fsm       <= FSM_WAIT_LOCK;
                ovrd      <= 1'd0;
                qpllreset <= 1'd1;
                qpllpd    <= 1'd0;
                end
            else
                begin
                fsm       <= FSM_IDLE;
                ovrd      <= ovrd;
                qpllreset <= &qpllreset_in_reg2;
                qpllpd    <= &qpllpd_in_reg2;
                end
            end  
            
        //---------- Wait for CPLL and QPLL to Lose Lock ---
        FSM_WAIT_LOCK :
        
            begin
            fsm       <= ((&(~cplllock_reg2)) && (&(~qplllock_reg2)) ? FSM_MMCM_LOCK : FSM_WAIT_LOCK);
            ovrd      <= ovrd;
            qpllreset <= qpllreset;
            qpllpd    <= qpllpd;
            end      
            
        //---------- Wait for MMCM and CPLL Lock -----------
        FSM_MMCM_LOCK :
        
            begin
            fsm       <= ((mmcm_lock_reg2 && (&cplllock_reg2)) ? FSM_DRP_START_NOM : FSM_MMCM_LOCK);
            ovrd      <= ovrd;
            qpllreset <= qpllreset;
            qpllpd    <= qpllpd;
            end      
            
        //---------- Start QPLL DRP for Normal QPLL Lock Mode 
        FSM_DRP_START_NOM:
        
            begin
            fsm       <= (&(~drp_done_reg2) ? FSM_DRP_DONE_NOM : FSM_DRP_START_NOM);
            ovrd      <= ovrd;
            qpllreset <= qpllreset;
            qpllpd    <= qpllpd;
            end

        //---------- Wait for QPLL DRP Done ----------------
        FSM_DRP_DONE_NOM :
        
            begin
            fsm       <= (&drp_done_reg2 ? FSM_QPLLLOCK : FSM_DRP_DONE_NOM);
            ovrd      <= ovrd;
            qpllreset <= qpllreset;
            qpllpd    <= qpllpd;
            end 
            
        //---------- Wait for QPLL Lock --------------------
        FSM_QPLLLOCK :
        
            begin
            fsm       <= (&qplllock_reg2 ? ((BYPASS_COARSE_OVRD == 1) ? FSM_QPLL_PDRESET : FSM_DRP_START_OPT) : FSM_QPLLLOCK);
            ovrd      <= ovrd;
            qpllreset <= 1'd0;
            qpllpd    <= qpllpd;
            end
            
        //---------- Start QPLL DRP for Optimized QPLL Lock Mode 
        FSM_DRP_START_OPT:
        
            begin
            fsm       <= (&(~drp_done_reg2) ? FSM_DRP_DONE_OPT : FSM_DRP_START_OPT);
            ovrd      <= 1'd1;
            qpllreset <= qpllreset;
            qpllpd    <= qpllpd;
            end

        //---------- Wait for QPLL DRP Done ----------------
        FSM_DRP_DONE_OPT :
        
            begin
            if (&drp_done_reg2)
                begin
                fsm       <= ((PCIE_PLL_SEL == "QPLL") ? FSM_QPLL_RESET : FSM_QPLL_PDRESET);
                ovrd      <= ovrd;
                qpllreset <= (PCIE_PLL_SEL == "QPLL");
                qpllpd    <= qpllpd;
                end
            else
                begin
                fsm       <= FSM_DRP_DONE_OPT;
                ovrd      <= ovrd;
                qpllreset <= qpllreset;
                qpllpd    <= qpllpd;
                end
            end 
            
        //---------- Reset QPLL ----------------------------
        FSM_QPLL_RESET :
            
            begin
            fsm       <= (&(~qplllock_reg2) ? FSM_QPLLLOCK2 : FSM_QPLL_RESET);  
            ovrd      <= ovrd;
            qpllreset <= 1'd1;
            qpllpd    <= 1'd0;
            end     
            
        //---------- Wait for QPLL Lock --------------------
        FSM_QPLLLOCK2 :
        
            begin
            fsm       <= (&qplllock_reg2 ? FSM_IDLE : FSM_QPLLLOCK2);
            ovrd      <= ovrd;
            qpllreset <= 1'd0;
            qpllpd    <= 1'd0;
            end
            
        //---------- Hold QPLL in Reset --------------------
        FSM_QPLL_PDRESET :
        
            begin
            fsm       <= FSM_QPLL_PD;
            ovrd      <= ovrd;
            qpllreset <= (PCIE_PLL_SEL == "CPLL") ? (rate_reg2 != 2'd2) : 1'd0; 
            qpllpd    <= qpllpd;
            end
            
        //---------- Power-down QPLL ----------------------- 
        FSM_QPLL_PD :
        
            begin
            fsm       <= FSM_IDLE;
            ovrd      <= ovrd;
            qpllreset <= qpllreset;
            qpllpd    <= (PCIE_PLL_SEL == "CPLL") ? (rate_reg2 != 2'd2) : 1'd0; 
            end 
                
        //---------- Default State -------------------------
        default :
        
            begin
            fsm       <= FSM_WAIT_LOCK;
            ovrd      <= 1'd0;
            qpllreset <= 1'd0;
            qpllpd    <= 1'd0;
            end

        endcase
        
        end
        
end



//---------- QPLL Lock Output --------------------------------------------------
assign QRST_OVRD          = ovrd;
assign QRST_DRP_START     = (fsm == FSM_DRP_START_NOM) || (fsm == FSM_DRP_START_OPT); 
assign QRST_QPLLRESET_OUT = qpllreset;
assign QRST_QPLLPD_OUT    = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : qpllpd);  
assign QRST_IDLE          = (fsm == FSM_IDLE);
assign QRST_FSM           = fsm;                   



endmodule



`timescale 1ns/1ps
module model_ap2_tst_pipe_user #
(

    parameter PCIE_SIM_MODE    = "FALSE",                   // PCIe sim mode 
    parameter PCIE_USE_MODE    = "3.0",                     // PCIe sim version
    parameter PCIE_OOBCLK_MODE = 1,                         // PCIe OOB clock mode
    parameter RXCDRLOCK_MAX    = 4'd15,                     // RXCDRLOCK max count
    parameter RXVALID_MAX      = 4'd15,                     // RXVALID max count
    parameter CONVERGE_MAX     = 22'd3125000                // Convergence max count
    
)

(

    //---------- Input -------------------------------------
    input               USER_TXUSRCLK,
    input               USER_RXUSRCLK,
    input               USER_OOBCLK_IN,
    input               USER_RST_N,
    input               USER_RXUSRCLK_RST_N,
    input               USER_PCLK_SEL,
    input               USER_RESETOVRD_START,
    input               USER_TXRESETDONE,
    input               USER_RXRESETDONE,
    input               USER_TXELECIDLE,
    input               USER_TXCOMPLIANCE,
    input               USER_RXCDRLOCK_IN,
    input               USER_RXVALID_IN,
    input               USER_RXSTATUS_IN,
    input               USER_PHYSTATUS_IN,
    input               USER_RATE_DONE, 
    input               USER_RST_IDLE,
    input               USER_RATE_RXSYNC,
    input               USER_RATE_IDLE,
    input               USER_RATE_GEN3,
    input               USER_RXEQ_ADAPT_DONE,
    
    //---------- Output ------------------------------------
    output              USER_OOBCLK,
    output              USER_RESETOVRD,
    output              USER_TXPMARESET,                            
    output              USER_RXPMARESET,                           
    output              USER_RXCDRRESET,               
    output              USER_RXCDRFREQRESET,           
    output              USER_RXDFELPMRESET,            
    output              USER_EYESCANRESET,             
    output              USER_TXPCSRESET,                              
    output              USER_RXPCSRESET,                            
    output              USER_RXBUFRESET,   
    output              USER_RESETOVRD_DONE,            
    output              USER_RESETDONE,
    output              USER_ACTIVE_LANE,
    output              USER_RXCDRLOCK_OUT,
    output              USER_RXVALID_OUT,
    output              USER_PHYSTATUS_OUT,
    output              USER_PHYSTATUS_RST,
    output              USER_GEN3_RDY,
    output              USER_RX_CONVERGE 

);
    
    //---------- Input Registers ---------------------------   
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 pclk_sel_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 resetovrd_start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxresetdone_reg1; 
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txelecidle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txcompliance_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxcdrlock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxvalid_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxstatus_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rst_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_rxsync_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_gen3_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_adapt_done_reg1;

(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 pclk_sel_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 resetovrd_start_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxresetdone_reg2; 
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txelecidle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txcompliance_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)	  reg	              rxcdrlock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxvalid_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxstatus_reg2; 
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_done_reg2;   
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rst_idle_reg2; 
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_rxsync_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_gen3_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_adapt_done_reg2;
    
    //---------- Internal Signal ---------------------------
    reg         [ 1:0]  oobclk_cnt    =  2'd0;
    reg         [ 7:0]  reset_cnt     =  8'd127;
    reg         [ 3:0]  rxcdrlock_cnt =  4'd0;
    reg         [ 3:0]  rxvalid_cnt   =  4'd0;
    reg         [21:0]  converge_cnt  = 22'd0;
    reg                 converge_gen3 =  1'd0;
    
    //---------- Output Registers --------------------------
    reg                 oobclk   = 1'd0;
    reg         [ 7:0]  reset    = 8'h00;
    reg                 gen3_rdy = 1'd0;
    reg         [ 1:0]  fsm      = 2'd0;
    
    //---------- FSM ---------------------------------------                                         
    localparam          FSM_IDLE       = 2'd0; 
    localparam          FSM_RESETOVRD  = 2'd1;
    localparam          FSM_RESET_INIT = 2'd2;
    localparam          FSM_RESET      = 2'd3;    
    
    //---------- Simulation Speedup ------------------------
    localparam converge_max_cnt = (PCIE_SIM_MODE == "TRUE") ? 22'd100 : CONVERGE_MAX;                                                              



//---------- Input FF ----------------------------------------------------------
always @ (posedge USER_TXUSRCLK)
begin

    if (!USER_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------  
        pclk_sel_reg1        <= 1'd0; 
        resetovrd_start_reg1 <= 1'd0;
        txresetdone_reg1     <= 1'd0;
        rxresetdone_reg1     <= 1'd0; 
        txelecidle_reg1      <= 1'd0;
        txcompliance_reg1    <= 1'd0;
        rxcdrlock_reg1 	     <= 1'd0;
        rxeq_adapt_done_reg1 <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        pclk_sel_reg2        <= 1'd0;
        resetovrd_start_reg2 <= 1'd0;
        txresetdone_reg2     <= 1'd0;
        rxresetdone_reg2     <= 1'd0; 
        txelecidle_reg2      <= 1'd0;
        txcompliance_reg2    <= 1'd0;
        rxcdrlock_reg2 	     <= 1'd0;
        rxeq_adapt_done_reg2 <= 1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        pclk_sel_reg1        <= USER_PCLK_SEL;
        resetovrd_start_reg1 <= USER_RESETOVRD_START;
        txresetdone_reg1     <= USER_TXRESETDONE;
        rxresetdone_reg1     <= USER_RXRESETDONE;
        txelecidle_reg1      <= USER_TXELECIDLE;
        txcompliance_reg1    <= USER_TXCOMPLIANCE;
        rxcdrlock_reg1 	     <= USER_RXCDRLOCK_IN;
        rxeq_adapt_done_reg1 <= USER_RXEQ_ADAPT_DONE;
        //---------- 2nd Stage FF --------------------------
        pclk_sel_reg2        <= pclk_sel_reg1;
        resetovrd_start_reg2 <= resetovrd_start_reg1;
        txresetdone_reg2     <= txresetdone_reg1;      
        rxresetdone_reg2     <= rxresetdone_reg1;      
        txelecidle_reg2      <= txelecidle_reg1;       
        txcompliance_reg2    <= txcompliance_reg1;  
        rxcdrlock_reg2 	     <= rxcdrlock_reg1;  
        rxeq_adapt_done_reg2 <= rxeq_adapt_done_reg1;
        end
        
end 



//---------- Input FF ----------------------------------------------------------
always @ (posedge USER_RXUSRCLK)
begin

    if (!USER_RXUSRCLK_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------   
        rxvalid_reg1     <= 1'd0;
        rxstatus_reg1    <= 1'd0;
        rst_idle_reg1    <= 1'd0; 
        rate_done_reg1   <= 1'd0;
        rate_rxsync_reg1 <= 1'd0;
        rate_idle_reg1   <= 1'd0;
        rate_gen3_reg1   <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        rxvalid_reg2     <= 1'd0;
        rxstatus_reg2    <= 1'd0;
        rst_idle_reg2    <= 1'd0; 
        rate_done_reg2   <= 1'd0;
        rate_rxsync_reg2 <= 1'd0;
        rate_idle_reg2   <= 1'd0;
        rate_gen3_reg2   <= 1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        rxvalid_reg1     <= USER_RXVALID_IN;
        rxstatus_reg1    <= USER_RXSTATUS_IN;
        rst_idle_reg1    <= USER_RST_IDLE; 
        rate_done_reg1   <= USER_RATE_DONE;
        rate_rxsync_reg1 <= USER_RATE_RXSYNC;
        rate_idle_reg1   <= USER_RATE_IDLE;
        rate_gen3_reg1   <= USER_RATE_GEN3;
        //---------- 2nd Stage FF --------------------------  	   
        rxvalid_reg2     <= rxvalid_reg1;            
        rxstatus_reg2    <= rxstatus_reg1; 
        rst_idle_reg2    <= rst_idle_reg1;
        rate_done_reg2   <= rate_done_reg1;  
        rate_rxsync_reg2 <= rate_rxsync_reg1;
        rate_idle_reg2   <= rate_idle_reg1;
        rate_gen3_reg2   <= rate_gen3_reg1;      
        end
        
end 



//---------- Generate Reset Override -------------------------------------------
generate if (PCIE_USE_MODE == "1.0") 

    begin : resetovrd

    //---------- Reset Counter -------------------------------------------------
    always @ (posedge USER_TXUSRCLK)
    begin
    
        if (!USER_RST_N)
            reset_cnt <= 8'd127;
        else
        
            //---------- Decrement Counter ---------------------
            if (((fsm == FSM_RESETOVRD) || (fsm == FSM_RESET)) && (reset_cnt != 8'd0))
                reset_cnt <= reset_cnt - 8'd1;
                
            //---------- Reset Counter -------------------------
            else 
            
                case (reset) 
                8'b00000000 : reset_cnt <= 8'd127;              // Programmable PMARESET       time
                8'b11111111 : reset_cnt <= 8'd127;              // Programmable RXCDRRESET     time
                8'b11111110 : reset_cnt <= 8'd127;              // Programmable RXCDRFREQRESET time
                8'b11111100 : reset_cnt <= 8'd127;              // Programmable RXDFELPMRESET  time
                8'b11111000 : reset_cnt <= 8'd127;              // Programmable EYESCANRESET   time
                8'b11110000 : reset_cnt <= 8'd127;              // Programmable PCSRESET       time
                8'b11100000 : reset_cnt <= 8'd127;              // Programmable RXBUFRESET     time
                8'b11000000 : reset_cnt <= 8'd127;              // Programmable RESETOVRD deassertion time
                8'b10000000 : reset_cnt <= 8'd127;
                default     : reset_cnt <= 8'd127; 
                endcase
                
    end 
    
    
    
    //---------- Reset Shift Register ------------------------------------------
    always @ (posedge USER_TXUSRCLK)
    begin
    
        if (!USER_RST_N)
            reset <= 8'h00;
        else
        
            //---------- Initialize Reset Register ---------
            if (fsm == FSM_RESET_INIT)
                reset <= 8'hFF;   
            //---------- Shift Reset Register --------------
            else if ((fsm == FSM_RESET) && (reset_cnt == 8'd0))
                reset <= {reset[6:0], 1'd0};        
            //---------- Hold Reset Register ---------------
            else
                reset <= reset;
            
    end
         
            
    
    //---------- Reset Override FSM --------------------------------------------
    always @ (posedge USER_TXUSRCLK)
    begin
    
        if (!USER_RST_N)
            fsm <= FSM_IDLE;     
                           
        else
        
            begin
            
            case (fsm)
            //---------- Idle State ------------------------
            FSM_IDLE       : fsm <= resetovrd_start_reg2 ? FSM_RESETOVRD : FSM_IDLE;
            //---------- Assert RESETOVRD ------------------
            FSM_RESETOVRD  : fsm <= (reset_cnt == 8'd0) ? FSM_RESET_INIT : FSM_RESETOVRD;
            //---------- Initialize Reset ------------------
            FSM_RESET_INIT : fsm <= FSM_RESET;
            //---------- Shift Reset -----------------------
            FSM_RESET      : fsm <= ((reset == 8'd0) && rxresetdone_reg2) ? FSM_IDLE : FSM_RESET;  
            //---------- Default State ---------------------
            default        : fsm <= FSM_IDLE;
        	  endcase
            
            end
    
    end
    
    end 

//---------- Disable Reset Override --------------------------------------------
else 

    begin : resetovrd_disble

    //---------- Generate Default Signals --------------------------------------
    always @ (posedge USER_TXUSRCLK)
    begin    
    
       if (!USER_RST_N)
           begin   
           reset_cnt <= 8'hFF;
           reset     <= 8'd0;
           fsm       <= 2'd0; 
           end
       else
           begin   
           reset_cnt <= 8'hFF;
           reset     <= 8'd0;
           fsm       <= 2'd0; 
           end
        
    end

    end

endgenerate



//---------- Generate OOB Clock Divider ------------------------
generate if (PCIE_OOBCLK_MODE == 1) 

    begin : oobclk_div
    
    //---------- OOB Clock Divider -----------------------------
    always @ (posedge USER_OOBCLK_IN)
    begin
    
        if (!USER_RST_N)
            begin
            oobclk_cnt <= 2'd0;
            oobclk     <= 1'd0;
            end
        else
            begin
            oobclk_cnt <= oobclk_cnt + 2'd1;
            oobclk     <= pclk_sel_reg2 ? oobclk_cnt[1] : oobclk_cnt[0];
            end
            
    end 
    
    end
   
else

    begin : oobclk_div_disable
    
    //---------- OOB Clock Default -------------------------
    always @ (posedge USER_OOBCLK_IN)
    begin
    
        if (!USER_RST_N)
            begin
            oobclk_cnt <= 2'd0;
            oobclk     <= 1'd0;
            end
        else
            begin
            oobclk_cnt <= 2'd0;
            oobclk     <= 1'd0;
            end
            
    end 
    
    end   
   
endgenerate

//---------- RXCDRLOCK Filter --------------------------------------------------
always @ (posedge USER_TXUSRCLK)
begin

    if (!USER_RST_N)
        rxcdrlock_cnt <= 4'd0;
    else
    
        //---------- Increment RXCDRLOCK Counter -----------
        if (rxcdrlock_reg2 && (rxcdrlock_cnt != RXCDRLOCK_MAX))
            rxcdrlock_cnt <= rxcdrlock_cnt + 4'd1;
            
        //---------- Hold RXCDRLOCK Counter ----------------
        else if (rxcdrlock_reg2 && (rxcdrlock_cnt == RXCDRLOCK_MAX))
            rxcdrlock_cnt <= rxcdrlock_cnt;
            
        //---------- Reset RXCDRLOCK Counter ---------------
        else
            rxcdrlock_cnt <= 4'd0;
        
end 



//---------- RXVALID Filter ----------------------------------------------------
always @ (posedge USER_RXUSRCLK)
begin

    if (!USER_RXUSRCLK_RST_N)
        rxvalid_cnt <= 4'd0;
    else
    
        //---------- Increment RXVALID Counter -------------
        if (rxvalid_reg2 && (rxvalid_cnt != RXVALID_MAX) && (!rxstatus_reg2))
            rxvalid_cnt <= rxvalid_cnt + 4'd1;
            
        //---------- Hold RXVALID Counter ------------------
        else if (rxvalid_reg2 && (rxvalid_cnt == RXVALID_MAX))
            rxvalid_cnt <= rxvalid_cnt;
            
        //---------- Reset RXVALID Counter -----------------
        else
            rxvalid_cnt <= 4'd0;
        
end 



//---------- Converge Counter --------------------------------------------------
always @ (posedge USER_TXUSRCLK)
begin

    if (!USER_RST_N)
        converge_cnt <= 22'd0;
    else
    
        //---------- Enter Gen1/Gen2 -----------------------
        if (rst_idle_reg2 && rate_idle_reg2 && !rate_gen3_reg2)
            begin
            
            //---------- Increment Converge Counter --------
            if (converge_cnt < converge_max_cnt) 
                converge_cnt <= converge_cnt + 22'd1;
            //---------- Hold Converge Counter -------------
            else 
                converge_cnt <= converge_cnt;
                
            end
            
        //---------- Reset Converge Counter ----------------
        else
            converge_cnt <= 22'd0;
        
end 



//---------- Converge ----------------------------------------------------------
always @ (posedge USER_TXUSRCLK)
begin

    if (!USER_RST_N)
        converge_gen3 <= 1'd0;
    else
    
        //---------- Enter Gen3 ----------------------------
        if (rate_gen3_reg2)
        
            //---------- Wait for RX equalization adapt done 
            if (rxeq_adapt_done_reg2)
                converge_gen3 <= 1'd1;
            else
                converge_gen3 <= converge_gen3;
        
        //-------- Exit Gen3 -------------------------------
        else
        
            converge_gen3 <= 1'd0;
        
        
end 



//---------- GEN3_RDY Generator ------------------------------------------------
always @ (posedge USER_RXUSRCLK)
begin

    if (!USER_RXUSRCLK_RST_N)
        gen3_rdy <= 1'd0;
    else   
        gen3_rdy <= rate_idle_reg2 && rate_gen3_reg2;    
        
end 



//---------- PIPE User Override Reset Output -----------------------------------  
assign USER_RESETOVRD      = (fsm != FSM_IDLE);
assign USER_TXPMARESET     = 1'd0; 
assign USER_RXPMARESET     = reset[0];  
assign USER_RXCDRRESET     = reset[1];
assign USER_RXCDRFREQRESET = reset[2];
assign USER_RXDFELPMRESET  = reset[3];
assign USER_EYESCANRESET   = reset[4];
assign USER_TXPCSRESET     = 1'd0;  
assign USER_RXPCSRESET     = reset[5];  
assign USER_RXBUFRESET     = reset[6];  
assign USER_RESETOVRD_DONE = (fsm == FSM_IDLE);

//---------- PIPE User Output --------------------------------------------------
assign USER_OOBCLK         = oobclk; 
assign USER_RESETDONE      = (txresetdone_reg2 && rxresetdone_reg2);
assign USER_ACTIVE_LANE    = !(txelecidle_reg2 && txcompliance_reg2);
//----------------------------------------------------------
assign USER_RXCDRLOCK_OUT  = (USER_RXCDRLOCK_IN && (rxcdrlock_cnt == RXCDRLOCK_MAX));        // Filtered RXCDRLOCK
//----------------------------------------------------------
assign USER_RXVALID_OUT    = ((USER_RXVALID_IN  && (rxvalid_cnt == RXVALID_MAX)) &&          // Filtered RXVALID
                              rst_idle_reg2                                      &&          // Force RXVALID = 0 during reset
                              rate_idle_reg2);                                               // Force RXVALID = 0 during rate change
//----------------------------------------------------------
assign USER_PHYSTATUS_OUT  = (!rst_idle_reg2                                              || // Force PHYSTATUS = 1 during reset
                              ((rate_idle_reg2 || rate_rxsync_reg2) && USER_PHYSTATUS_IN) || // Raw PHYSTATUS
                              rate_done_reg2);                                               // Gated PHYSTATUS for rate change
//----------------------------------------------------------
assign USER_PHYSTATUS_RST  = !rst_idle_reg2;                                                 // Filtered PHYSTATUS for reset
//----------------------------------------------------------
assign USER_GEN3_RDY       = 0;//gen3_rdy;                                                      
//----------------------------------------------------------
assign USER_RX_CONVERGE    = (converge_cnt == converge_max_cnt) || converge_gen3;   



endmodule


`timescale 1ns/1ps
module model_ap2_tst_gtp_pipe_rate #
(

    parameter PCIE_SIM_SPEEDUP = "FALSE",                   // PCIe sim mode 
    parameter TXDATA_WAIT_MAX  = 4'd15                      // TXDATA wait max

)

(

    //---------- Input -------------------------------------
    input               RATE_CLK,
    input               RATE_RST_N,
    input       [ 1:0]  RATE_RATE_IN,
    input               RATE_DRP_DONE,
    input               RATE_RXPMARESETDONE,
    input               RATE_TXRATEDONE,
    input               RATE_RXRATEDONE,
    input               RATE_TXSYNC_DONE,
    input               RATE_PHYSTATUS,
    
    //---------- Output ------------------------------------
    output              RATE_PCLK_SEL,
    output              RATE_DRP_START,
    output              RATE_DRP_X16,
    output      [ 2:0]  RATE_RATE_OUT,
    output              RATE_TXSYNC_START,
    output              RATE_DONE,
    output              RATE_IDLE,
    output      [ 4:0]  RATE_FSM

);

    //---------- Input FF or Buffer ------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_in_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 drp_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxpmaresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txratedone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxratedone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 phystatus_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_done_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_in_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 drp_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxpmaresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txratedone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxratedone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 phystatus_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_done_reg2;
    
    //---------- Internal Signals --------------------------
    wire        [ 2:0]  rate;
    reg         [ 3:0]  txdata_wait_cnt = 4'd0;
    reg                 txratedone      = 1'd0;
    reg                 rxratedone      = 1'd0;
    reg                 phystatus       = 1'd0;
    reg                 ratedone        = 1'd0;
    
    //---------- Output FF or Buffer -----------------------
    reg                 pclk_sel =  1'd0; 
    reg         [ 2:0]  rate_out =  3'd0; 
    reg         [ 3:0]  fsm      =  0;                 
   
    //---------- FSM ---------------------------------------                                         
    localparam          FSM_IDLE           = 0; 
    localparam          FSM_TXDATA_WAIT    = 1;           
    localparam          FSM_PCLK_SEL       = 2; 
    localparam          FSM_DRP_X16_START  = 3;
    localparam          FSM_DRP_X16_DONE   = 4;   
    localparam          FSM_RATE_SEL       = 5;
    localparam          FSM_RXPMARESETDONE = 6; 
    localparam          FSM_DRP_X20_START  = 7;
    localparam          FSM_DRP_X20_DONE   = 8;   
    localparam          FSM_RATE_DONE      = 9;
    localparam          FSM_TXSYNC_START   = 10;
    localparam          FSM_TXSYNC_DONE    = 11;             
    localparam          FSM_DONE           = 12; // Must sync value to pipe_user.v
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin    
        //---------- 1st Stage FF -------------------------- 
        rate_in_reg1        <= 2'd0;
        drp_done_reg1       <= 1'd0;
        rxpmaresetdone_reg1 <= 1'd0;
        txratedone_reg1     <= 1'd0;
        rxratedone_reg1     <= 1'd0;
        phystatus_reg1      <= 1'd0;
        txsync_done_reg1    <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        rate_in_reg2        <= 2'd0;
        drp_done_reg2       <= 1'd0;
        rxpmaresetdone_reg2 <= 1'd0;
        txratedone_reg2     <= 1'd0;
        rxratedone_reg2     <= 1'd0;
        phystatus_reg2      <= 1'd0;
        txsync_done_reg2    <= 1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        rate_in_reg1        <= RATE_RATE_IN;
        drp_done_reg1       <= RATE_DRP_DONE;
        rxpmaresetdone_reg1 <= RATE_RXPMARESETDONE;
        txratedone_reg1     <= RATE_TXRATEDONE;
        rxratedone_reg1     <= RATE_RXRATEDONE;
        phystatus_reg1      <= RATE_PHYSTATUS;
        txsync_done_reg1    <= RATE_TXSYNC_DONE;
        //---------- 2nd Stage FF --------------------------
        rate_in_reg2        <= rate_in_reg1;
        drp_done_reg2       <= drp_done_reg1;
        rxpmaresetdone_reg2 <= rxpmaresetdone_reg1;
        txratedone_reg2     <= txratedone_reg1;
        rxratedone_reg2     <= rxratedone_reg1;
        phystatus_reg2      <= phystatus_reg1;
        txsync_done_reg2    <= txsync_done_reg1;   
        end
        
end    



//---------- Select Rate -------------------------------------------------------
//  Gen1 :  div 2 using [TX/RX]OUT_DIV = 2
//  Gen2 :  div 1 using [TX/RX]RATE = 3'd1
//------------------------------------------------------------------------------
assign rate = (rate_in_reg2 == 2'd1) ? 3'd1 : 3'd0;



//---------- TXDATA Wait Counter -----------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        txdata_wait_cnt <= 4'd0;
    else
    
        //---------- Increment Wait Counter ----------------
        if ((fsm == FSM_TXDATA_WAIT) && (txdata_wait_cnt < TXDATA_WAIT_MAX))
            txdata_wait_cnt <= txdata_wait_cnt + 4'd1;
            
        //---------- Hold Wait Counter ---------------------
        else if ((fsm == FSM_TXDATA_WAIT) && (txdata_wait_cnt == TXDATA_WAIT_MAX))
            txdata_wait_cnt <= txdata_wait_cnt;
            
        //---------- Reset Wait Counter --------------------
        else
            txdata_wait_cnt <= 4'd0;
        
end 



//---------- Latch TXRATEDONE, RXRATEDONE, and PHYSTATUS -----------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin   
        txratedone <= 1'd0;
        rxratedone <= 1'd0; 
        phystatus  <= 1'd0;
        ratedone   <= 1'd0;
        end
    else
        begin  

        if ((fsm == FSM_RATE_DONE) || (fsm == FSM_RXPMARESETDONE) || (fsm == FSM_DRP_X20_START) || (fsm == FSM_DRP_X20_DONE))
        
            begin
            
            //---------- Latch TXRATEDONE ------------------
            if (txratedone_reg2)
                txratedone <= 1'd1; 
            else
                txratedone <= txratedone;
 
            //---------- Latch RXRATEDONE ------------------
            if (rxratedone_reg2)
                rxratedone <= 1'd1; 
            else
                rxratedone <= rxratedone;
  
            //---------- Latch PHYSTATUS -------------------
            if (phystatus_reg2)
                phystatus <= 1'd1; 
            else
                phystatus <= phystatus;
  
            //---------- Latch Rate Done -------------------
            if (rxratedone && txratedone && phystatus)
                ratedone <= 1'd1; 
            else
                ratedone <= ratedone;
  
            end
  
        else 
        
            begin
            txratedone <= 1'd0;
            rxratedone <= 1'd0;
            phystatus  <= 1'd0;
            ratedone   <= 1'd0;
            end
        
        end
        
end    



//---------- PIPE Rate FSM -----------------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin
        fsm      <= FSM_IDLE;
        pclk_sel <= 1'd0; 
        rate_out <= 3'd0;                              
        end
    else
        begin
        
        case (fsm)
            
        //---------- Idle State ----------------------------
        FSM_IDLE :
        
            begin
            //---------- Detect Rate Change ----------------
            if (rate_in_reg2 != rate_in_reg1)
                begin
                fsm      <= FSM_TXDATA_WAIT;
                pclk_sel <= pclk_sel;
                rate_out <= rate_out;
                end
            else
                begin
                fsm      <= FSM_IDLE;
                pclk_sel <= pclk_sel;
                rate_out <= rate_out;
                end
            end 
            
        //---------- Wait for TXDATA to TX[P/N] Latency ----    
        FSM_TXDATA_WAIT :
        
            begin
            fsm      <= (txdata_wait_cnt == TXDATA_WAIT_MAX) ? FSM_PCLK_SEL : FSM_TXDATA_WAIT;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end 

        //---------- Select PCLK Frequency -----------------
        //  Gen1 : PCLK = 125 MHz
        //  Gen2 : PCLK = 250 MHz
        //--------------------------------------------------
        FSM_PCLK_SEL :
        
            begin
            fsm      <= (PCIE_SIM_SPEEDUP == "TRUE") ? FSM_RATE_SEL : FSM_DRP_X16_START;    
            pclk_sel <= (rate_in_reg2 == 2'd1);
            rate_out <= rate_out;
            end
            
        //---------- Start DRP x16 -------------------------
        FSM_DRP_X16_START :
            
            begin
            fsm      <= (!drp_done_reg2) ? FSM_DRP_X16_DONE : FSM_DRP_X16_START;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end
            
        //---------- Wait for DRP x16 Done -----------------    
        FSM_DRP_X16_DONE :
        
            begin  
            fsm      <= drp_done_reg2 ? FSM_RATE_SEL : FSM_DRP_X16_DONE;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end      

        //---------- Select Rate ---------------------------
        FSM_RATE_SEL :
        
            begin
            fsm      <= (PCIE_SIM_SPEEDUP == "TRUE") ? FSM_RATE_DONE : FSM_RXPMARESETDONE;
            pclk_sel <= pclk_sel;
            rate_out <= rate;                               // Update [TX/RX]RATE
            end    
            
        //---------- Wait for RXPMARESETDONE De-assertion --
        FSM_RXPMARESETDONE :
        
            begin
            fsm      <= (!rxpmaresetdone_reg2) ? FSM_DRP_X20_START : FSM_RXPMARESETDONE;  
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end  
            
        //---------- Start DRP x20 -------------------------
        FSM_DRP_X20_START :
            
            begin
            fsm      <= (!drp_done_reg2) ? FSM_DRP_X20_DONE : FSM_DRP_X20_START;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end
            
        //---------- Wait for DRP x20 Done -----------------    
        FSM_DRP_X20_DONE :
        
            begin  
            fsm      <= drp_done_reg2 ? FSM_RATE_DONE : FSM_DRP_X20_DONE;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end      
            
        //---------- Wait for Rate Change Done ------------- 
        FSM_RATE_DONE :
        
            begin
            if (ratedone) 
                fsm <= FSM_TXSYNC_START;
            else      
                fsm <= FSM_RATE_DONE;
            
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end      
            
        //---------- Start TX Sync -------------------------
        FSM_TXSYNC_START:
        
            begin
            fsm      <= (!txsync_done_reg2 ? FSM_TXSYNC_DONE : FSM_TXSYNC_START);
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end
            
        //---------- Wait for TX Sync Done -----------------
        FSM_TXSYNC_DONE:
        
            begin
            fsm      <= (txsync_done_reg2 ? FSM_DONE : FSM_TXSYNC_DONE);
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end        

        //---------- Rate Change Done ----------------------
        FSM_DONE :  
          
            begin  
            fsm      <= FSM_IDLE;
            pclk_sel <= pclk_sel;
            rate_out <= rate_out;
            end
               
        //---------- Default State -------------------------
        default :
        
            begin
            fsm      <= FSM_IDLE;
            pclk_sel <= 1'd0; 
            rate_out <= 3'd0;  
            end

        endcase
        
        end
        
end 



//---------- PIPE Rate Output --------------------------------------------------
assign RATE_PCLK_SEL     = pclk_sel;
assign RATE_DRP_START    = (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X20_START); 
assign RATE_DRP_X16      = (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X16_DONE);
assign RATE_RATE_OUT     = rate_out;
assign RATE_TXSYNC_START = (fsm == FSM_TXSYNC_START);
assign RATE_DONE         = (fsm == FSM_DONE);
assign RATE_IDLE         = (fsm == FSM_IDLE);
assign RATE_FSM          = {1'd0, fsm};   



endmodule



`timescale 1ns/1ps
module model_ap2_tst_pipe_rate #
(

    parameter PCIE_SIM_SPEEDUP  = "FALSE",                  // PCIe sim speedup
    parameter PCIE_GT_DEVICE    = "GTX",                    // PCIe GT device
    parameter PCIE_USE_MODE     = "3.0",                    // PCIe use mode
    parameter PCIE_PLL_SEL      = "CPLL",                   // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_POWER_SAVING = "TRUE",                   // PCIe power saving
    parameter PCIE_ASYNC_EN     = "FALSE",                  // PCIe async enable
    parameter PCIE_TXBUF_EN     = "FALSE",                  // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_RXBUF_EN     = "TRUE",                   // PCIe RX buffer enable for Gen3      only
    parameter TXDATA_WAIT_MAX   = 4'd15                     // TXDATA wait max

)

(

    //---------- Input -------------------------------------
    input               RATE_CLK,
    input               RATE_RST_N,
    input               RATE_RST_IDLE,
    input               RATE_ACTIVE_LANE,
    input       [ 1:0]  RATE_RATE_IN,
    input               RATE_CPLLLOCK,
    input               RATE_QPLLLOCK,
    input               RATE_MMCM_LOCK,
    input               RATE_DRP_DONE,
    input               RATE_RXPMARESETDONE,
    input               RATE_TXRESETDONE,
    input               RATE_RXRESETDONE,
    input               RATE_TXRATEDONE,
    input               RATE_RXRATEDONE,
    input               RATE_PHYSTATUS,
    input               RATE_RESETOVRD_DONE,
    input               RATE_TXSYNC_DONE,
    input               RATE_RXSYNC_DONE,
    
    //---------- Output ------------------------------------
    output              RATE_CPLLPD,
    output              RATE_QPLLPD,
    output              RATE_CPLLRESET,
    output              RATE_QPLLRESET,
    output              RATE_TXPMARESET,
    output              RATE_RXPMARESET,
    output              RATE_DRP_START,
    output      [ 1:0]  RATE_SYSCLKSEL,
    output              RATE_PCLK_SEL,
    output              RATE_GEN3,
    output              RATE_DRP_X16X20_MODE,
    output              RATE_DRP_X16,
    output      [ 2:0]  RATE_RATE_OUT,
    output              RATE_RESETOVRD_START,
    output              RATE_TXSYNC_START,
    output              RATE_DONE,
    output              RATE_RXSYNC_START,
    output              RATE_RXSYNC,
    output              RATE_IDLE,
    output      [ 4:0]  RATE_FSM

);

    //---------- Input FF or Buffer ------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rst_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_in_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 cplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 qplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 mmcm_lock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 drp_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxpmaresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txratedone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxratedone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 phystatus_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 resetovrd_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_done_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsync_done_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rst_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_in_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 cplllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 qplllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 mmcm_lock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 drp_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxpmaresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txratedone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxratedone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 phystatus_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 resetovrd_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_done_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsync_done_reg2;
    
    //---------- Internal Signals --------------------------
    wire                pll_lock;
    wire        [ 2:0]  rate;
    reg         [ 3:0]  txdata_wait_cnt = 4'd0;
    reg                 txratedone      = 1'd0;
    reg                 rxratedone      = 1'd0;
    reg                 phystatus       = 1'd0;
    reg                 ratedone        = 1'd0;
    reg                 gen3_exit       = 1'd0;
    
    //---------- Output FF or Buffer -----------------------
    reg                 cpllpd     =  1'd0;
    reg                 qpllpd     =  1'd0;
    reg                 cpllreset  =  1'd0;
    reg                 qpllreset  =  1'd0;
    reg                 txpmareset =  1'd0;
    reg                 rxpmareset =  1'd0;
    reg         [ 1:0]  sysclksel  = (PCIE_PLL_SEL == "QPLL") ? 2'd1 : 2'd0;  
    reg                 gen3       =  1'd0;
    reg                 pclk_sel   =  1'd0; 
    reg         [ 2:0]  rate_out   =  3'd0; 
    reg                 drp_start       = 1'd0;
    reg                 drp_x16x20_mode = 1'd0;
    reg                 drp_x16         = 1'd0;
    reg         [4:0]   fsm             = 0;                 
   
    //---------- FSM ---------------------------------------        
    localparam          FSM_IDLE               = 0;
    localparam          FSM_PLL_PU             = 1; // Gen 3 only
    localparam          FSM_PLL_PURESET        = 2; // Gen 3 only
    localparam          FSM_PLL_LOCK           = 3; // Gen 3 or reset only
    localparam          FSM_DRP_X16_GEN3_START = 4;
    localparam          FSM_DRP_X16_GEN3_DONE  = 5;
    localparam          FSM_PMARESET_HOLD      = 6; // Gen 3 or reset only
    localparam          FSM_PLL_SEL            = 7; // Gen 3 or reset only
    localparam          FSM_MMCM_LOCK          = 8; // Gen 3 or reset only
    localparam          FSM_DRP_START          = 9; // Gen 3 or reset only
    localparam          FSM_DRP_DONE           = 10; // Gen 3 or reset only
    localparam          FSM_PMARESET_RELEASE   = 11; // Gen 3 only
    localparam          FSM_PMARESET_DONE      = 12; // Gen 3 only
    localparam          FSM_TXDATA_WAIT        = 13;
    localparam          FSM_PCLK_SEL           = 14;
    localparam          FSM_DRP_X16_START      = 15;
    localparam          FSM_DRP_X16_DONE       = 16;
    localparam          FSM_RATE_SEL           = 17;
    localparam          FSM_RXPMARESETDONE     = 18;
    localparam          FSM_DRP_X20_START      = 19;
    localparam          FSM_DRP_X20_DONE       = 20;
    localparam          FSM_RATE_DONE          = 21;
    localparam          FSM_RESETOVRD_START    = 22; // PCIe use mode 1.0 only
    localparam          FSM_RESETOVRD_DONE     = 23; // PCIe use mode 1.0 only
    localparam          FSM_PLL_PDRESET        = 24;
    localparam          FSM_PLL_PD             = 25;
    localparam          FSM_TXSYNC_START       = 26;
    localparam          FSM_TXSYNC_DONE        = 27;
    localparam          FSM_DONE               = 28; // Must sync value to pipe_user.v
    localparam          FSM_RXSYNC_START       = 29; // Gen 3 only
    localparam          FSM_RXSYNC_DONE        = 30; // Gen 3 only                                 
    
    
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin    
        //---------- 1st Stage FF -------------------------- 
        rst_idle_reg1       <= 1'd0;   
        rate_in_reg1        <= 2'd0;
        cplllock_reg1       <= 1'd0;
        qplllock_reg1       <= 1'd0;
        mmcm_lock_reg1      <= 1'd0;
        drp_done_reg1       <= 1'd0;
        rxpmaresetdone_reg1 <= 1'd0;
        txresetdone_reg1    <= 1'd0;
        rxresetdone_reg1    <= 1'd0;
        txratedone_reg1     <= 1'd0;
        rxratedone_reg1     <= 1'd0;
        phystatus_reg1      <= 1'd0;
        resetovrd_done_reg1 <= 1'd0; 
        txsync_done_reg1    <= 1'd0;
        rxsync_done_reg1    <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        rst_idle_reg2       <= 1'd0;
        rate_in_reg2        <= 2'd0;
        cplllock_reg2       <= 1'd0;
        qplllock_reg2       <= 1'd0;
        mmcm_lock_reg2      <= 1'd0;
        drp_done_reg2       <= 1'd0;
        rxpmaresetdone_reg2 <= 1'd0;
        txresetdone_reg2    <= 1'd0;
        rxresetdone_reg2    <= 1'd0;
        txratedone_reg2     <= 1'd0;
        rxratedone_reg2     <= 1'd0;
        phystatus_reg2      <= 1'd0;
        resetovrd_done_reg2 <= 1'd0;
        txsync_done_reg2    <= 1'd0;
        rxsync_done_reg2    <= 1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        rst_idle_reg1       <= RATE_RST_IDLE;
        rate_in_reg1        <= RATE_RATE_IN;
        cplllock_reg1       <= RATE_CPLLLOCK;
        qplllock_reg1       <= RATE_QPLLLOCK;
        mmcm_lock_reg1      <= RATE_MMCM_LOCK;
        drp_done_reg1       <= RATE_DRP_DONE;
        rxpmaresetdone_reg1 <= RATE_RXPMARESETDONE;
        txresetdone_reg1    <= RATE_TXRESETDONE;
        rxresetdone_reg1    <= RATE_RXRESETDONE;
        txratedone_reg1     <= RATE_TXRATEDONE;
        rxratedone_reg1     <= RATE_RXRATEDONE;
        phystatus_reg1      <= RATE_PHYSTATUS;
        resetovrd_done_reg1 <= RATE_RESETOVRD_DONE;
        txsync_done_reg1    <= RATE_TXSYNC_DONE;
        rxsync_done_reg1    <= RATE_RXSYNC_DONE;
        //---------- 2nd Stage FF --------------------------
        rst_idle_reg2       <= rst_idle_reg1;
        rate_in_reg2        <= rate_in_reg1;
        cplllock_reg2       <= cplllock_reg1;
        qplllock_reg2       <= qplllock_reg1;
        mmcm_lock_reg2      <= mmcm_lock_reg1;
        drp_done_reg2       <= drp_done_reg1;
        rxpmaresetdone_reg2 <= rxpmaresetdone_reg1;
        txresetdone_reg2    <= txresetdone_reg1;
        rxresetdone_reg2    <= rxresetdone_reg1;
        txratedone_reg2     <= txratedone_reg1;
        rxratedone_reg2     <= rxratedone_reg1;
        phystatus_reg2      <= phystatus_reg1;
        resetovrd_done_reg2 <= resetovrd_done_reg1;
        txsync_done_reg2    <= txsync_done_reg1;   
        rxsync_done_reg2    <= rxsync_done_reg1; 
        end
        
end    



//---------- Select CPLL or QPLL Lock ------------------------------------------
//  Gen1 : Wait for QPLL lock if QPLL is used for Gen1/Gen2, else wait for CPLL lock 
//  Gen2 : Wait for QPLL lock if QPLL is used for Gen1/Gen2, else wait for CPLL lock
//  Gen3 : Wait for QPLL lock
//------------------------------------------------------------------------------
assign pll_lock = (rate_in_reg2 == 2'd2) || (PCIE_PLL_SEL == "QPLL") ? qplllock_reg2 : cplllock_reg2;



//---------- Select Rate -------------------------------------------------------
//  Gen1 : Div 4 using [TX/RX]OUT_DIV = 4 if QPLL is used for Gen1/Gen2, else div 2 using [TX/RX]OUT_DIV = 2
//  Gen2 : Div 2 using [TX/RX]RATE = 3'd2 if QPLL is used for Gen1/Gen2, else div 1 using [TX/RX]RATE = 3'd1
//  Gen3 : Div 1 using [TX/RX]OUT_DIV = 1
//------------------------------------------------------------------------------
assign rate = (rate_in_reg2 == 2'd1) && (PCIE_PLL_SEL == "QPLL") ? 3'd2 : 
              (rate_in_reg2 == 2'd1) && (PCIE_PLL_SEL == "CPLL") ? 3'd1 : 3'd0;



//---------- TXDATA Wait Counter -----------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        txdata_wait_cnt <= 4'd0;
    else
    
        //---------- Increment Wait Counter ----------------
        if ((fsm == FSM_TXDATA_WAIT) && (txdata_wait_cnt < TXDATA_WAIT_MAX))
            txdata_wait_cnt <= txdata_wait_cnt + 4'd1;
            
        //---------- Hold Wait Counter ---------------------
        else if ((fsm == FSM_TXDATA_WAIT) && (txdata_wait_cnt == TXDATA_WAIT_MAX))
            txdata_wait_cnt <= txdata_wait_cnt;
            
        //---------- Reset Wait Counter --------------------
        else
            txdata_wait_cnt <= 4'd0;
        
end 



//---------- Latch TXRATEDONE, RXRATEDONE, and PHYSTATUS -----------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin   
        txratedone <= 1'd0;
        rxratedone <= 1'd0; 
        phystatus  <= 1'd0;
        ratedone   <= 1'd0;
        end
    else
        begin  

        if (fsm == FSM_RATE_DONE)
        
            begin
            
            //---------- Latch TXRATEDONE ------------------
            if (txratedone_reg2)
                txratedone <= 1'd1; 
            else
                txratedone <= txratedone;
 
            //---------- Latch RXRATEDONE ------------------
            if (rxratedone_reg2)
                rxratedone <= 1'd1; 
            else
                rxratedone <= rxratedone;
  
            //---------- Latch PHYSTATUS -------------------
            if (phystatus_reg2)
                phystatus <= 1'd1; 
            else
                phystatus <= phystatus;
  
            //---------- Latch Rate Done -------------------
            if (rxratedone && txratedone && phystatus)
                ratedone <= 1'd1; 
            else
                ratedone <= ratedone;
  
            end
  
        else 
        
            begin
            txratedone <= 1'd0;
            rxratedone <= 1'd0;
            phystatus  <= 1'd0;
            ratedone   <= 1'd0;
            end
        
        end
        
end    



//---------- PIPE Rate FSM -----------------------------------------------------
always @ (posedge RATE_CLK)
begin

    if (!RATE_RST_N)
        begin
        fsm        <= FSM_PLL_LOCK;
        gen3_exit  <= 1'd0;
        cpllpd     <= 1'd0;
        qpllpd     <= 1'd0;
        cpllreset  <= 1'd0;
        qpllreset  <= 1'd0;
        txpmareset <= 1'd0;
        rxpmareset <= 1'd0;
        sysclksel  <= (PCIE_PLL_SEL == "QPLL") ? 2'd1 : 2'd0;                               
        pclk_sel   <= 1'd0; 
        gen3       <= 1'd0;
        rate_out   <= 3'd0;  
        drp_start       <= 1'd0;
        drp_x16x20_mode <= 1'd0;  
        drp_x16         <= 1'd0;                          
        end
    else
        begin
        
        case (fsm)
            
        //---------- Idle State ----------------------------
        FSM_IDLE :
        
            begin
            //---------- Detect Rate Change ----------------
            if (rate_in_reg2 != rate_in_reg1)
                begin
                fsm        <= ((rate_in_reg2 == 2'd2) || (rate_in_reg1 == 2'd2)) ? FSM_PLL_PU : FSM_TXDATA_WAIT;
                gen3_exit  <= (rate_in_reg2 == 2'd2); 
                cpllpd     <= cpllpd;
                qpllpd     <= qpllpd;
                cpllreset  <= cpllreset;
                qpllreset  <= qpllreset;
                txpmareset <= txpmareset;
                rxpmareset <= rxpmareset;
                sysclksel  <= sysclksel;
                pclk_sel   <= pclk_sel;
                gen3       <= gen3;
                rate_out   <= rate_out;
                drp_start       <= 1'd0;
                drp_x16x20_mode <= 1'd0;
                drp_x16         <= 1'd0;    
                end
            else
                begin
                fsm        <= FSM_IDLE;
                gen3_exit  <= gen3_exit;
                cpllpd     <= cpllpd;
                qpllpd     <= qpllpd;
                cpllreset  <= cpllreset;
                qpllreset  <= qpllreset;
                txpmareset <= txpmareset;
                rxpmareset <= rxpmareset;
                sysclksel  <= sysclksel;
                pclk_sel   <= pclk_sel;
                gen3       <= gen3;
                rate_out   <= rate_out;
                drp_start       <= 1'd0;
                drp_x16x20_mode <= 1'd0;
                drp_x16         <= 1'd0;    
                end
            end 
            
        //---------- Power-up PLL --------------------------
        FSM_PLL_PU :
        
            begin
            fsm        <= FSM_PLL_PURESET;
            gen3_exit  <= gen3_exit;
            cpllpd     <= (PCIE_PLL_SEL == "QPLL");
            qpllpd     <= 1'd0;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end  
            
        //---------- Release PLL Resets --------------------
        FSM_PLL_PURESET :
        
            begin
            fsm        <= FSM_PLL_LOCK;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= (PCIE_PLL_SEL == "QPLL");
            qpllreset  <= 1'd0;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end 

        //---------- Wait for PLL Lock ---------------------
        FSM_PLL_LOCK :
        
            begin
            fsm        <= (pll_lock ? ((!rst_idle_reg2 || (rate_in_reg2 == 2'd1)) ? FSM_PMARESET_HOLD : FSM_DRP_X16_GEN3_START) : FSM_PLL_LOCK);  
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Start DRP x16 -------------------------
        FSM_DRP_X16_GEN3_START :
            
            begin
            fsm        <= (!drp_done_reg2) ? FSM_DRP_X16_GEN3_DONE : FSM_DRP_X16_GEN3_START;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd1;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd1;    
            end
            
        //---------- Wait for DRP x16 Done -----------------    
        FSM_DRP_X16_GEN3_DONE :
        
            begin  
            fsm        <= drp_done_reg2 ? FSM_PMARESET_HOLD : FSM_DRP_X16_GEN3_DONE;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd1;    
            end  

        //---------- Hold both PMA in Reset ----------------
        //  Gen1 : Release PMA Reset
        //  Gen2 : Release PMA Reset
        //  Gen3 : Hold PMA Reset
        //--------------------------------------------------
        FSM_PMARESET_HOLD :
        
            begin
            fsm        <= FSM_PLL_SEL;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= ((rate_in_reg2 == 2'd2) || gen3_exit);
            rxpmareset <= ((rate_in_reg2 == 2'd2) || gen3_exit);
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Select PLL ----------------------------
        //  Gen1 : QPLL if PCIE_PLL_SEL = QPLL, else CPLL
        //  Gen2 : QPLL if PCIE_PLL_SEL = QPLL, else CPLL
        //  Gen3 : QPLL
        //--------------------------------------------------
        FSM_PLL_SEL :
        
            begin
            fsm        <= FSM_MMCM_LOCK;    
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= ((rate_in_reg2 == 2'd2) || (PCIE_PLL_SEL == "QPLL")) ? 2'd1 : 2'd0;                          
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Check for MMCM Lock -------------------
        FSM_MMCM_LOCK :
        
            begin
            fsm        <= (mmcm_lock_reg2 && !rxpmaresetdone_reg2 ? FSM_DRP_START : FSM_MMCM_LOCK);  
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Start DRP -----------------------------
        FSM_DRP_START:
        
            begin
            fsm        <= (!drp_done_reg2 ? FSM_DRP_DONE : FSM_DRP_START);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= ((rate_in_reg2 == 2'd1) || (rate_in_reg2 == 2'd2));
            gen3       <= (rate_in_reg2 == 2'd2);  
            rate_out   <= (((rate_in_reg2 == 2'd2) || gen3_exit) ? rate : rate_out);  
            drp_start       <= 1'd1;
            drp_x16x20_mode <= 1'd0;  
            drp_x16         <= 1'd0;                     
            end

        //---------- Wait for DRP Done ---------------------
        FSM_DRP_DONE :
        
            begin
            fsm        <= ((drp_done_reg2 && pll_lock) ? (rst_idle_reg2 ? FSM_PMARESET_RELEASE : FSM_IDLE): FSM_DRP_DONE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end 

        //---------- Release PMA Resets --------------------
        FSM_PMARESET_RELEASE :
        
            begin
            fsm        <= FSM_PMARESET_DONE;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= 1'd0;
            rxpmareset <= 1'd0;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Wait for both TX/RX PMA Reset Dones and PHYSTATUS Deassertion
        FSM_PMARESET_DONE :
        
            begin
            fsm        <= (((rxresetdone_reg2 && txresetdone_reg2 && !phystatus_reg2) || !RATE_ACTIVE_LANE) ? FSM_TXDATA_WAIT : FSM_PMARESET_DONE); 
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Wait for TXDATA to TX[P/N] Latency ----
        FSM_TXDATA_WAIT :
        
            begin
            fsm        <= (txdata_wait_cnt == TXDATA_WAIT_MAX) ? FSM_PCLK_SEL : FSM_TXDATA_WAIT;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end 

        //---------- Select PCLK Frequency -----------------
        //  Gen1 : PCLK = 125 MHz
        //  Gen2 : PCLK = 250 MHz
        //  Gen3 : PCLK = 250 MHz
        //--------------------------------------------------
        FSM_PCLK_SEL :
        
            begin
            fsm        <= ((PCIE_GT_DEVICE == "GTH") && ((rate_in_reg2 == 2'd1) || ((!gen3_exit) && (rate_in_reg2 == 2'd0)))) ? FSM_DRP_X16_START : FSM_RATE_SEL; 
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= ((rate_in_reg2 == 2'd1) || (rate_in_reg2 == 2'd2));
            gen3       <= gen3;    
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;    
            end

        //---------- Start DRP x16 -------------------------
        FSM_DRP_X16_START :
            
            begin
            fsm        <= (!drp_done_reg2) ? FSM_DRP_X16_DONE : FSM_DRP_X16_START;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd1;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd1;
            end
            
        //---------- Wait for DRP x16 Done -----------------    
        FSM_DRP_X16_DONE :
        
            begin  
            fsm        <= drp_done_reg2 ? FSM_RATE_SEL : FSM_DRP_X16_DONE;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd1;
            end    

        //---------- Select Rate ---------------------------
        FSM_RATE_SEL :
        
            begin
            fsm        <= ((PCIE_GT_DEVICE == "GTH") && ((rate_in_reg2 == 2'd1) || ((!gen3_exit) && (rate_in_reg2 == 2'd0)))) ? FSM_RXPMARESETDONE : FSM_RATE_DONE;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate;                             // Update [TX/RX]RATE
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end    
            
        //---------- Wait for RXPMARESETDONE De-assertion --
        FSM_RXPMARESETDONE :
        
            begin
            fsm        <= (!rxpmaresetdone_reg2) ? FSM_DRP_X20_START : FSM_RXPMARESETDONE;  
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end  
            
        //---------- Start DRP x20 -------------------------
        FSM_DRP_X20_START :
            
            begin
            fsm        <= (!drp_done_reg2) ? FSM_DRP_X20_DONE : FSM_DRP_X20_START;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd1;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd0;
            end
            
        //---------- Wait for DRP x20 Done -----------------    
        FSM_DRP_X20_DONE :
        
            begin  
            fsm        <= drp_done_reg2 ? FSM_RATE_DONE : FSM_DRP_X20_DONE;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd1;
            drp_x16         <= 1'd0;
            end       
            
        //---------- Wait for Rate Change Done ------------- 
        FSM_RATE_DONE :
        
            begin
            if (ratedone || (rate_in_reg2 == 2'd2) || (gen3_exit) || !RATE_ACTIVE_LANE) 
                if ((PCIE_USE_MODE == "1.0") && (rate_in_reg2 != 2'd2) && (!gen3_exit)) 
                    fsm <= FSM_RESETOVRD_START;
                else
                    fsm <= FSM_PLL_PDRESET;  
            else      
                fsm <= FSM_RATE_DONE;
            
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end      
            
        //---------- Reset Override Start ------------------
        FSM_RESETOVRD_START:
        
            begin
            fsm        <= (!resetovrd_done_reg2 ? FSM_RESETOVRD_DONE : FSM_RESETOVRD_START);    
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end
            
        //---------- Reset Override Done -------------------
        FSM_RESETOVRD_DONE :
        
            begin
            fsm        <= (resetovrd_done_reg2 ? FSM_PLL_PDRESET : FSM_RESETOVRD_DONE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end  
                
        //---------- Hold PLL Not Used in Reset ------------
        FSM_PLL_PDRESET :
        
            begin
            fsm        <= FSM_PLL_PD;
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= (PCIE_PLL_SEL == "QPLL") ? 1'd1 : (rate_in_reg2 == 2'd2);
            qpllreset  <= (PCIE_PLL_SEL == "QPLL") ? 1'd0 : (rate_in_reg2 != 2'd2);
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end    
            
        //---------- Power-Down PLL Not Used ---------------
        FSM_PLL_PD :
        
            begin
            fsm        <= (((rate_in_reg2 == 2'd2) || (PCIE_TXBUF_EN == "FALSE")) ? FSM_TXSYNC_START : FSM_DONE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= (PCIE_PLL_SEL == "QPLL") ? 1'd1 : (rate_in_reg2 == 2'd2);
            qpllpd     <= (PCIE_PLL_SEL == "QPLL") ? 1'd0 : (rate_in_reg2 != 2'd2);
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end         
            
        //---------- Start TX Sync -------------------------
        FSM_TXSYNC_START:
        
            begin
            fsm        <= (!txsync_done_reg2 ? FSM_TXSYNC_DONE : FSM_TXSYNC_START);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end
            
        //---------- Wait for TX Sync Done -----------------
        FSM_TXSYNC_DONE:
        
            begin
            fsm        <= (txsync_done_reg2 ? FSM_DONE : FSM_TXSYNC_DONE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end        

        //---------- Rate Change Done ----------------------
        FSM_DONE :  
          
            begin  
            fsm        <= (((rate_in_reg2 == 2'd2) && (PCIE_RXBUF_EN == "FALSE") && (PCIE_ASYNC_EN == "TRUE")) ? FSM_RXSYNC_START : FSM_IDLE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end
               
        //---------- Start RX Sync -------------------------
        FSM_RXSYNC_START:
        
            begin
            fsm        <= (!rxsync_done_reg2 ? FSM_RXSYNC_DONE : FSM_RXSYNC_START);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end
            
        //---------- Wait for RX Sync Done -----------------
        FSM_RXSYNC_DONE:
        
            begin          
            fsm        <= (rxsync_done_reg2 ? FSM_IDLE : FSM_RXSYNC_DONE);
            gen3_exit  <= gen3_exit;
            cpllpd     <= cpllpd;
            qpllpd     <= qpllpd;
            cpllreset  <= cpllreset;
            qpllreset  <= qpllreset;
            txpmareset <= txpmareset;
            rxpmareset <= rxpmareset;
            sysclksel  <= sysclksel;
            pclk_sel   <= pclk_sel;
            gen3       <= gen3;
            rate_out   <= rate_out;
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end   
                
        //---------- Default State -------------------------
        default :
        
            begin
            fsm        <= FSM_IDLE;
            gen3_exit  <= 1'd0;
            cpllpd     <= 1'd0;
            qpllpd     <= 1'd0;
            cpllreset  <= 1'd0;
            qpllreset  <= 1'd0;
            txpmareset <= 1'd0;
            rxpmareset <= 1'd0;
            sysclksel  <= (PCIE_PLL_SEL == "QPLL") ? 2'd1 : 2'd0;                               
            pclk_sel   <= 1'd0; 
            gen3       <= 1'd0;
            rate_out   <= 3'd0;  
            drp_start       <= 1'd0;
            drp_x16x20_mode <= 1'd0;
            drp_x16         <= 1'd0;
            end

        endcase
        
        end
        
end 



//---------- PIPE Rate Output --------------------------------------------------
assign RATE_CPLLPD          = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : cpllpd);
assign RATE_QPLLPD          = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : qpllpd);
assign RATE_CPLLRESET       = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : cpllreset);
assign RATE_QPLLRESET       = ((PCIE_POWER_SAVING == "FALSE") ? 1'd0 : qpllreset);
assign RATE_TXPMARESET      = txpmareset;
assign RATE_RXPMARESET      = rxpmareset;
assign RATE_SYSCLKSEL       = sysclksel;

//assign RATE_DRP_START       = (fsm == FSM_DRP_START) || (fsm == FSM_DRP_X16_GEN3_START) || (fsm == FSM_DRP_X16_START) || (fsm == FSM_DRP_X20_START); 
  assign RATE_DRP_START       = drp_start;

//assign RATE_DRP_X16X20_MODE = (fsm == FSM_DRP_X16_GEN3_START) || (fsm == FSM_DRP_X16_GEN3_DONE) ||
//                              (fsm == FSM_DRP_X16_START)      || (fsm == FSM_DRP_X16_DONE) || 
//                              (fsm == FSM_DRP_X20_START)      || (fsm == FSM_DRP_X20_DONE);
  assign RATE_DRP_X16X20_MODE = drp_x16x20_mode;

//assign RATE_DRP_X16         = (fsm == FSM_DRP_X16_GEN3_START) || (fsm == FSM_DRP_X16_GEN3_DONE) ||
//                              (fsm == FSM_DRP_X16_START)      || (fsm == FSM_DRP_X16_DONE);
  assign RATE_DRP_X16         = drp_x16;  
                          
assign RATE_PCLK_SEL        = pclk_sel;
assign RATE_GEN3            = gen3;
assign RATE_RATE_OUT        = rate_out;
assign RATE_RESETOVRD_START = (fsm == FSM_RESETOVRD_START);
assign RATE_TXSYNC_START    = (fsm == FSM_TXSYNC_START);
assign RATE_DONE            = (fsm == FSM_DONE);
assign RATE_RXSYNC_START    = (fsm == FSM_RXSYNC_START);
assign RATE_RXSYNC          = ((fsm == FSM_RXSYNC_START) || (fsm == FSM_RXSYNC_DONE));
assign RATE_IDLE            = (fsm == FSM_IDLE);
assign RATE_FSM             = fsm;   



endmodule


`timescale 1ns/1ps
module model_ap2_tst_pipe_sync #
(

    parameter PCIE_GT_DEVICE       = "GTX",                 // PCIe GT device
    parameter PCIE_TXBUF_EN        = "FALSE",               // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_RXBUF_EN        = "TRUE",                // PCIe TX buffer enable for Gen3      only
    parameter PCIE_TXSYNC_MODE     = 0,                     // PCIe TX sync mode
    parameter PCIE_RXSYNC_MODE     = 0,                     // PCIe RX sync mode
    parameter PCIE_LANE            = 1,                     // PCIe lane
    parameter PCIE_LINK_SPEED      = 3,                     // PCIe link speed
    parameter BYPASS_TXDELAY_ALIGN = 0,                     // Bypass TX delay align
    parameter BYPASS_RXDELAY_ALIGN = 0                      // Bypass RX delay align

)

(

    //---------- Input -------------------------------------
    input               SYNC_CLK,
    input               SYNC_RST_N,
    input               SYNC_SLAVE,
    input               SYNC_GEN3,
    input               SYNC_RATE_IDLE,
    input               SYNC_MMCM_LOCK,
    input               SYNC_RXELECIDLE,
    input               SYNC_RXCDRLOCK,
    input               SYNC_ACTIVE_LANE,
    
    input               SYNC_TXSYNC_START,
    input               SYNC_TXPHINITDONE,   
    input               SYNC_TXDLYSRESETDONE,
    input               SYNC_TXPHALIGNDONE,
    input               SYNC_TXSYNCDONE,
        
    input               SYNC_RXSYNC_START,
    input               SYNC_RXDLYSRESETDONE,
    input               SYNC_RXPHALIGNDONE_M,
    input               SYNC_RXPHALIGNDONE_S,
    input               SYNC_RXSYNC_DONEM_IN,
    input               SYNC_RXSYNCDONE,
    
    //---------- Output ------------------------------------
    output              SYNC_TXPHDLYRESET,
    output              SYNC_TXPHALIGN,     
    output              SYNC_TXPHALIGNEN,  
    output              SYNC_TXPHINIT,       
    output              SYNC_TXDLYBYPASS,  
    output              SYNC_TXDLYSRESET,
    output              SYNC_TXDLYEN,   
    output              SYNC_TXSYNC_DONE,
    output    [ 5:0]    SYNC_FSM_TX,
    
    output              SYNC_RXPHALIGN,
    output              SYNC_RXPHALIGNEN,
    output              SYNC_RXDLYBYPASS,
    output              SYNC_RXDLYSRESET,
    output              SYNC_RXDLYEN,
    output              SYNC_RXDDIEN,
    output              SYNC_RXSYNC_DONEM_OUT,
    output              SYNC_RXSYNC_DONE,
    output    [ 6:0]    SYNC_FSM_RX

);          

    //---------- Input Register ----------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_idle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg		      mmcm_lock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxelecidle_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxcdrlock_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg2;     
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rate_idle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg		      mmcm_lock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxelecidle_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxcdrlock_reg2;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg		      txsync_start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphinitdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txdlysresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphaligndone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsyncdone_reg1;
                                                   
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_start_reg2;     
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphinitdone_reg2;     
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txdlysresetdone_reg2;    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphaligndone_reg2;   
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsyncdone_reg2; 
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsync_start_reg3;     
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphinitdone_reg3;     
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txdlysresetdone_reg3;    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txphaligndone_reg3;   
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 txsyncdone_reg3;     
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg		      rxsync_start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxdlysresetdone_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxphaligndone_m_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxphaligndone_s_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsync_donem_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsyncdone_reg1;

(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg		      rxsync_start_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxdlysresetdone_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxphaligndone_m_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxphaligndone_s_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsync_donem_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxsyncdone_reg2;
    
    //---------- Output Register ---------------------------          
    reg                 txdlyen     = 1'd0;
    reg                 txsync_done = 1'd0;
    reg         [ 5:0]  fsm_tx      = 6'd0;     
    
    reg                 rxdlyen     = 1'd0;
    reg                 rxsync_done = 1'd0;         
    reg	        [ 6:0]  fsm_rx      = 7'd0;   
   
    //---------- FSM ---------------------------------------                                         
    localparam          FSM_TXSYNC_IDLE  = 6'b000001; 
    localparam          FSM_MMCM_LOCK    = 6'b000010;                                     
    localparam          FSM_TXSYNC_START = 6'b000100;
    localparam          FSM_TXPHINITDONE = 6'b001000;       // Manual TX sync only
    localparam          FSM_TXSYNC_DONE1 = 6'b010000;   
    localparam          FSM_TXSYNC_DONE2 = 6'b100000;             
        
    localparam          FSM_RXSYNC_IDLE  = 7'b0000001; 
    localparam          FSM_RXCDRLOCK    = 7'b0000010;                                     
    localparam          FSM_RXSYNC_START = 7'b0000100;
    localparam          FSM_RXSYNC_DONE1 = 7'b0001000;                                     
    localparam          FSM_RXSYNC_DONE2 = 7'b0010000;
    localparam          FSM_RXSYNC_DONES = 7'b0100000;
    localparam          FSM_RXSYNC_DONEM = 7'b1000000;
        
    
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge SYNC_CLK)
begin

    if (!SYNC_RST_N)
        begin    
        //---------- 1st Stage FF --------------------------  
        gen3_reg1            <= 1'd0;
        rate_idle_reg1       <= 1'd0;
        mmcm_lock_reg1       <= 1'd0;
        rxelecidle_reg1      <= 1'd0;
        rxcdrlock_reg1 	     <= 1'd0;
 
        txsync_start_reg1	   <= 1'd0;
        txphinitdone_reg1    <= 1'd0;
        txdlysresetdone_reg1 <= 1'd0;
        txphaligndone_reg1   <= 1'd0;
        txsyncdone_reg1      <= 1'd0;
        
        rxsync_start_reg1	   <= 1'd0; 
        rxdlysresetdone_reg1 <= 1'd0;
        rxphaligndone_m_reg1 <= 1'd0;
        rxphaligndone_s_reg1 <= 1'd0;
        rxsync_donem_reg1    <= 1'd0;    
        rxsyncdone_reg1      <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        gen3_reg2            <= 1'd0;
        rate_idle_reg2       <= 1'd0;
        mmcm_lock_reg2       <= 1'd0;
        rxelecidle_reg2      <= 1'd0;
        rxcdrlock_reg2 	     <= 1'd0;
        
        txsync_start_reg2	   <= 1'd0;
        txphinitdone_reg2    <= 1'd0;
        txdlysresetdone_reg2 <= 1'd0;
        txphaligndone_reg2   <= 1'd0;
        txsyncdone_reg2      <= 1'd0;
        
        rxsync_start_reg2	   <= 1'd0; 
        rxdlysresetdone_reg2 <= 1'd0;
        rxphaligndone_m_reg2 <= 1'd0;
        rxphaligndone_s_reg2 <= 1'd0;
        rxsync_donem_reg2    <= 1'd0;
        rxsyncdone_reg2      <= 1'd0;
        //---------- 3rd Stage FF --------------------------
        txsync_start_reg3	   <= 1'd0;
        txphinitdone_reg3    <= 1'd0;
        txdlysresetdone_reg3 <= 1'd0;
        txphaligndone_reg3   <= 1'd0;
        txsyncdone_reg3      <= 1'd0;
        
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        gen3_reg1            <= SYNC_GEN3;
        rate_idle_reg1       <= SYNC_RATE_IDLE;
        mmcm_lock_reg1       <= SYNC_MMCM_LOCK;
        rxelecidle_reg1      <= SYNC_RXELECIDLE; 
        rxcdrlock_reg1       <= SYNC_RXCDRLOCK;

        txsync_start_reg1    <= SYNC_TXSYNC_START;
        txphinitdone_reg1    <= SYNC_TXPHINITDONE;
        txdlysresetdone_reg1 <= SYNC_TXDLYSRESETDONE;
        txphaligndone_reg1   <= SYNC_TXPHALIGNDONE;
        txsyncdone_reg1      <= SYNC_TXSYNCDONE;
        
        rxsync_start_reg1	   <= SYNC_RXSYNC_START; 
        rxdlysresetdone_reg1 <= SYNC_RXDLYSRESETDONE;
        rxphaligndone_m_reg1 <= SYNC_RXPHALIGNDONE_M;
        rxphaligndone_s_reg1 <= SYNC_RXPHALIGNDONE_S;
        rxsync_donem_reg1    <= SYNC_RXSYNC_DONEM_IN;
        rxsyncdone_reg1      <= SYNC_RXSYNCDONE; 
        //---------- 2nd Stage FF --------------------------
        gen3_reg2            <= gen3_reg1;
        rate_idle_reg2       <= rate_idle_reg1;
        mmcm_lock_reg2       <= mmcm_lock_reg1;
        rxelecidle_reg2      <= rxelecidle_reg1;
        rxcdrlock_reg2       <= rxcdrlock_reg1;
        
        txsync_start_reg2    <= txsync_start_reg1;       
        txphinitdone_reg2    <= txphinitdone_reg1; 
        txdlysresetdone_reg2 <= txdlysresetdone_reg1;   
        txphaligndone_reg2   <= txphaligndone_reg1;
        txsyncdone_reg2      <= txsyncdone_reg1;
        
        rxsync_start_reg2    <= rxsync_start_reg1;
        rxdlysresetdone_reg2 <= rxdlysresetdone_reg1; 
        rxphaligndone_m_reg2 <= rxphaligndone_m_reg1;
        rxphaligndone_s_reg2 <= rxphaligndone_s_reg1;
        rxsync_donem_reg2    <= rxsync_donem_reg1; 
        rxsyncdone_reg2      <= rxsyncdone_reg1;
        //---------- 3rd Stage FF --------------------------
        txsync_start_reg3    <= txsync_start_reg2;	   
        txphinitdone_reg3    <= txphinitdone_reg2;    
        txdlysresetdone_reg3 <= txdlysresetdone_reg2; 
        txphaligndone_reg3   <= txphaligndone_reg2;   
        txsyncdone_reg3      <= txsyncdone_reg2;      
        end
        
end       



//---------- Generate TX Sync FSM ----------------------------------------------
generate if ((PCIE_LINK_SPEED == 3) || (PCIE_TXBUF_EN == "FALSE")) 

    begin : txsync_fsm

    //---------- PIPE TX Sync FSM ----------------------------------------------
    always @ (posedge SYNC_CLK)
    begin
    
        if (!SYNC_RST_N)
            begin
            fsm_tx      <= FSM_TXSYNC_IDLE;   
            txdlyen     <= 1'd0; 
            txsync_done <= 1'd0;
            end                    
        else
            begin
            
            case (fsm_tx)
            
            //---------- Idle State ------------------------
            FSM_TXSYNC_IDLE :
            
                begin     
                //---------- Exiting Reset or Rate Change --
                if (txsync_start_reg2)
                    begin
                    fsm_tx      <= FSM_MMCM_LOCK;
                    txdlyen     <= 1'd0; 
                    txsync_done <= 1'd0;
                    end
                else
                    begin
                    fsm_tx      <= FSM_TXSYNC_IDLE;
                    txdlyen     <= txdlyen; 
                    txsync_done <= txsync_done;
                    end
                end
                
            //---------- Check MMCM Lock -------------------
            FSM_MMCM_LOCK :
            
                begin
                fsm_tx      <= (mmcm_lock_reg2 ? FSM_TXSYNC_START : FSM_MMCM_LOCK);
                txdlyen     <= 1'd0; 
                txsync_done <= 1'd0;  
                end
                
            //---------- TX Delay Soft Reset --------------- 
            FSM_TXSYNC_START :
            
                begin
                fsm_tx      <= (((!txdlysresetdone_reg3 && txdlysresetdone_reg2) || (((PCIE_GT_DEVICE == "GTH") || (PCIE_GT_DEVICE == "GTP")) && (PCIE_TXSYNC_MODE == 1) && SYNC_SLAVE)) ? FSM_TXPHINITDONE : FSM_TXSYNC_START);
                txdlyen     <= 1'd0; 
                txsync_done <= 1'd0;
                end
                
            //---------- Wait for TX Phase Init Done (Manual Mode Only)
            FSM_TXPHINITDONE :
            
                begin
                fsm_tx      <= (((!txphinitdone_reg3 && txphinitdone_reg2) || (PCIE_TXSYNC_MODE == 1) || (!SYNC_ACTIVE_LANE)) ? FSM_TXSYNC_DONE1 : FSM_TXPHINITDONE);
                txdlyen     <= 1'd0; 
                txsync_done <= 1'd0;
                end
                
            //---------- Wait for TX Phase Alignment Done --
            FSM_TXSYNC_DONE1 :
            
                begin
                if (((PCIE_GT_DEVICE == "GTH") || (PCIE_GT_DEVICE == "GTP")) && (PCIE_TXSYNC_MODE == 1) && !SYNC_SLAVE)
                   fsm_tx <= ((!txsyncdone_reg3 && txsyncdone_reg2)       || (!SYNC_ACTIVE_LANE) ? FSM_TXSYNC_DONE2 : FSM_TXSYNC_DONE1); 
                else
                   fsm_tx <= ((!txphaligndone_reg3 && txphaligndone_reg2) || (!SYNC_ACTIVE_LANE) ? FSM_TXSYNC_DONE2 : FSM_TXSYNC_DONE1); 
                
                txdlyen     <= 1'd0; 
                txsync_done <= 1'd0;
                end  
                
            //---------- Wait for Master TX Delay Alignment Done 
            FSM_TXSYNC_DONE2 :
            
                begin
                if ((!txphaligndone_reg3 && txphaligndone_reg2) || (!SYNC_ACTIVE_LANE) || SYNC_SLAVE || (((PCIE_GT_DEVICE == "GTH") || (PCIE_GT_DEVICE == "GTP")) && (PCIE_TXSYNC_MODE == 1)) || (BYPASS_TXDELAY_ALIGN == 1)) 
                    begin
                    fsm_tx      <= FSM_TXSYNC_IDLE;
                    txdlyen     <= !SYNC_SLAVE; 
                    txsync_done <= 1'd1;
                    end
                else
                    begin
                    fsm_tx      <= FSM_TXSYNC_DONE2;
                    txdlyen     <= !SYNC_SLAVE; 
                    txsync_done <= 1'd0;
                    end
                end         
                              
            //---------- Default State ---------------------
            default :
                begin 
                fsm_tx      <= FSM_TXSYNC_IDLE;
                txdlyen     <= 1'd0; 
                txsync_done <= 1'd0;
                end
                
            endcase
            
            end
            
    end     

    end  
          
//---------- TX Sync FSM Default------------------------------------------------
else 

    begin : txsync_fsm_disable
       
    //---------- Default -------------------------------------------------------
    always @ (posedge SYNC_CLK)
    begin    
        fsm_tx      <= FSM_TXSYNC_IDLE;
        txdlyen     <= 1'd0;
        txsync_done <= 1'd0; 
    end

    end 

endgenerate  

          
       
//---------- Generate RX Sync FSM ----------------------------------------------
generate if ((PCIE_LINK_SPEED == 3) && (PCIE_RXBUF_EN == "FALSE")) 

    begin : rxsync_fsm
   
    //---------- PIPE RX Sync FSM ----------------------------------------------
    always @ (posedge SYNC_CLK)
    begin
    
        if (!SYNC_RST_N)
            begin
            fsm_rx      <= FSM_RXSYNC_IDLE; 
            rxdlyen     <= 1'd0;
            rxsync_done <= 1'd0;   
            end                    
        else
            begin
            
            case (fsm_rx)
            
            //---------- Idle State ------------------------
            FSM_RXSYNC_IDLE :
            
                begin
                //---------- Exiting Rate Change -----------
                if (rxsync_start_reg2)
                    begin
                    fsm_rx      <= FSM_RXCDRLOCK;
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd0;
                    end
                //---------- Exiting Electrical Idle without Rate Change 
                else if (gen3_reg2 && rate_idle_reg2 && ((rxelecidle_reg2 == 1'd1) && (rxelecidle_reg1 == 1'd0)))
                    begin
                    fsm_rx      <= FSM_RXCDRLOCK;
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd0;   
                    end 
                //---------- Idle --------------------------
                else                    
                    begin
                    fsm_rx      <= FSM_RXSYNC_IDLE;
                    rxdlyen     <= rxelecidle_reg2 ? 1'd0 : rxdlyen;
                    rxsync_done <= rxelecidle_reg2 ? 1'd0 : rxsync_done;
                    end
                end
                
            //---------- Wait for RX Electrical Idle Exit and RX CDR Lock 
            FSM_RXCDRLOCK :
            
                begin
                fsm_rx      <= ((!rxelecidle_reg2 && rxcdrlock_reg2) ? FSM_RXSYNC_START : FSM_RXCDRLOCK);
                rxdlyen     <= 1'd0;
                rxsync_done <= 1'd0;
                end
                
            //---------- Start RX Sync with RX Delay Soft Reset
            FSM_RXSYNC_START :
            
                begin
                fsm_rx      <= ((!rxdlysresetdone_reg2 && rxdlysresetdone_reg1) ? FSM_RXSYNC_DONE1 : FSM_RXSYNC_START);
                rxdlyen     <= 1'd0;
                rxsync_done <= 1'd0;
                end     
                      
            //---------- Wait for RX Phase Alignment Done --
            FSM_RXSYNC_DONE1 :
            
                begin
                if (SYNC_SLAVE)
                    begin
                    fsm_rx      <= ((!rxphaligndone_s_reg2 && rxphaligndone_s_reg1) ? FSM_RXSYNC_DONE2 : FSM_RXSYNC_DONE1);
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd0;
                    end
                else
                    begin
                    fsm_rx      <= ((!rxphaligndone_m_reg2 && rxphaligndone_m_reg1) ? FSM_RXSYNC_DONE2 : FSM_RXSYNC_DONE1);
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd0;
                    end
                end  
                
            //---------- Wait for Master RX Delay Alignment Done 
            FSM_RXSYNC_DONE2 :
            
                begin   
                if (SYNC_SLAVE)
                    begin
                    fsm_rx      <= FSM_RXSYNC_IDLE;
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd1;
                    end
                else if ((!rxphaligndone_m_reg2 && rxphaligndone_m_reg1) || (BYPASS_RXDELAY_ALIGN == 1)) 
                    begin
                    fsm_rx      <= ((PCIE_LANE == 1) ? FSM_RXSYNC_IDLE : FSM_RXSYNC_DONES);
                    rxdlyen     <=  (PCIE_LANE == 1);
                    rxsync_done <=  (PCIE_LANE == 1);
                    end
                else
                    begin
                    fsm_rx      <= FSM_RXSYNC_DONE2;
                    rxdlyen     <= 1'd1;
                    rxsync_done <= 1'd0;
                    end
                end     
                
            //---------- Wait for Slave RX Phase Alignment Done 
            FSM_RXSYNC_DONES :
            
                begin
                if (!rxphaligndone_s_reg2 && rxphaligndone_s_reg1) 
                    begin
                    fsm_rx      <= FSM_RXSYNC_DONEM;
                    rxdlyen     <= 1'd1;
                    rxsync_done <= 1'd0;
                    end
                else
                    begin
                    fsm_rx      <= FSM_RXSYNC_DONES;
                    rxdlyen     <= 1'd0;
                    rxsync_done <= 1'd0;
                    end
                end           
                   
            //---------- Wait for Master RX Delay Alignment Done 
            FSM_RXSYNC_DONEM :
            
                begin
                if ((!rxphaligndone_m_reg2 && rxphaligndone_m_reg1) || (BYPASS_RXDELAY_ALIGN == 1)) 
                    begin
                    fsm_rx      <= FSM_RXSYNC_IDLE;
                    rxdlyen     <= 1'd1;
                    rxsync_done <= 1'd1;
                    end
                else
                    begin
                    fsm_rx      <= FSM_RXSYNC_DONEM;
                    rxdlyen     <= 1'd1;
                    rxsync_done <= 1'd0;
                    end
                end         
                              
            //---------- Default State ---------------------
            default : 
                begin
                fsm_rx      <= FSM_RXSYNC_IDLE;
                rxdlyen     <= 1'd0;
                rxsync_done <= 1'd0;
                end    
                        
        	   endcase
            
            end
            
    end            
        
    end  
          
//---------- RX Sync FSM Default -----------------------------------------------
else 

    begin : rxsync_fsm_disable
       
    //---------- Default -------------------------------------------------------
    always @ (posedge SYNC_CLK)
    begin    
        fsm_rx      <= FSM_RXSYNC_IDLE;
        rxdlyen     <= 1'd0;
        rxsync_done <= 1'd0; 
    end

    end 

endgenerate      
   


//---------- PIPE Sync Output --------------------------------------------------            
assign SYNC_TXPHALIGNEN      = ((PCIE_TXSYNC_MODE == 1) || (!gen3_reg2 && (PCIE_TXBUF_EN == "TRUE"))) ? 1'd0 : 1'd1;   
assign SYNC_TXDLYBYPASS      = 1'd0;                     
//assign SYNC_TXDLYSRESET    = !(((PCIE_GT_DEVICE == "GTH") || (PCIE_GT_DEVICE == "GTP")) && (PCIE_TXSYNC_MODE == 1) && SYNC_SLAVE) ? (fsm_tx == FSM_TXSYNC_START) : 1'd0; 
assign SYNC_TXDLYSRESET      = (fsm_tx == FSM_TXSYNC_START);
assign SYNC_TXPHDLYRESET     =  (((PCIE_GT_DEVICE == "GTH") || (PCIE_GT_DEVICE == "GTP")) && (PCIE_TXSYNC_MODE == 1) && SYNC_SLAVE) ? (fsm_tx == FSM_TXSYNC_START) : 1'd0;   
assign SYNC_TXPHINIT         = PCIE_TXSYNC_MODE ? 1'd0 : (fsm_tx == FSM_TXPHINITDONE); 
assign SYNC_TXPHALIGN        = PCIE_TXSYNC_MODE ? 1'd0 : (fsm_tx == FSM_TXSYNC_DONE1);
assign SYNC_TXDLYEN          = PCIE_TXSYNC_MODE ? 1'd0 : txdlyen;
assign SYNC_TXSYNC_DONE      = txsync_done;
assign SYNC_FSM_TX           = fsm_tx;

assign SYNC_RXPHALIGNEN      = ((PCIE_RXSYNC_MODE == 1) || (!gen3_reg2) || (PCIE_RXBUF_EN == "TRUE")) ? 1'd0 : 1'd1;  
assign SYNC_RXDLYBYPASS      = !gen3_reg2 || (PCIE_RXBUF_EN == "TRUE");
assign SYNC_RXDLYSRESET      = (fsm_rx == FSM_RXSYNC_START);
assign SYNC_RXPHALIGN        = PCIE_RXSYNC_MODE ? 1'd0 : (!SYNC_SLAVE ? (fsm_rx == FSM_RXSYNC_DONE1) : (rxsync_donem_reg2 && (fsm_rx == FSM_RXSYNC_DONE1)));
assign SYNC_RXDLYEN          = PCIE_RXSYNC_MODE ? 1'd0 : rxdlyen;
assign SYNC_RXDDIEN          = gen3_reg2 && (PCIE_RXBUF_EN == "FALSE"); 
assign SYNC_RXSYNC_DONE      = rxsync_done;
assign SYNC_RXSYNC_DONEM_OUT = (fsm_rx == FSM_RXSYNC_DONES);
assign SYNC_FSM_RX	         = fsm_rx;  



endmodule



`timescale 1ns/1ps
module model_ap2_tst_gtp_pipe_drp #
(

    parameter LOAD_CNT_MAX     = 2'd1,                      // Load max count
    parameter INDEX_MAX        = 1'd0                       // Index max count
    
)

(
    
    //---------- Input -------------------------------------
    input               DRP_CLK,
    input               DRP_RST_N,
    input               DRP_X16,
    input               DRP_START,
    input       [15:0]  DRP_DO,
    input               DRP_RDY,
    
    //---------- Output ------------------------------------
    output      [ 8:0]  DRP_ADDR,
    output              DRP_EN,  
    output      [15:0]  DRP_DI,   
    output              DRP_WE,
    output              DRP_DONE,
    output      [ 2:0]  DRP_FSM
    
);

    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg2;
    
    //---------- Internal Signals --------------------------
    reg         [ 1:0]  load_cnt =  2'd0;
    reg         [ 4:0]  index    =  5'd0;
    reg         [ 8:0]  addr_reg =  9'd0;
    reg         [15:0]  di_reg   = 16'd0;
    
    //---------- Output Registers --------------------------
    reg                 done     =  1'd0;
    reg         [ 2:0]  fsm      =  0;      
                        
    //---------- DRP Address -------------------------------          
    localparam          ADDR_RX_DATAWIDTH  = 9'h011;              
    
    //---------- DRP Mask ----------------------------------
    localparam          MASK_RX_DATAWIDTH  = 16'b1111011111111111;  // Unmask bit [   11]  
         
    //---------- DRP Data for x16 --------------------------
    localparam          X16_RX_DATAWIDTH   = 16'b0000000000000000;  // 2-byte (16-bit) internal data width
    
    //---------- DRP Data for x20 --------------------------                                  
    localparam          X20_RX_DATAWIDTH   = 16'b0000100000000000;  // 2-byte (20-bit) internal data width               
      
    //---------- DRP Data ----------------------------------                  
    wire        [15:0]  data_rx_datawidth;                 
           
    //---------- FSM ---------------------------------------  
    localparam          FSM_IDLE  = 0;  
    localparam          FSM_LOAD  = 1;                           
    localparam          FSM_READ  = 2;
    localparam          FSM_RRDY  = 3;
    localparam          FSM_WRITE = 4;
    localparam          FSM_WRDY  = 5;    
    localparam          FSM_DONE  = 6;   

    
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        //---------- 1st Stage FF --------------------------
        x16_reg1   <=  1'd0;
        do_reg1    <= 16'd0;
        rdy_reg1   <=  1'd0;
        start_reg1 <=  1'd0;
        //---------- 2nd Stage FF --------------------------
        x16_reg2   <=  1'd0;
        do_reg2    <= 16'd0;
        rdy_reg2   <=  1'd0;
        start_reg2 <=  1'd0;
        end
        
    else
        begin
        //---------- 1st Stage FF --------------------------
        x16_reg1   <= DRP_X16;
        do_reg1    <= DRP_DO;
        rdy_reg1   <= DRP_RDY;
        start_reg1 <= DRP_START;
        //---------- 2nd Stage FF --------------------------
        x16_reg2   <= x16_reg1;
        do_reg2    <= do_reg1;
        rdy_reg2   <= rdy_reg1;
        start_reg2 <= start_reg1;
        end
    
end  



//---------- Select DRP Data ---------------------------------------------------
assign data_rx_datawidth = x16_reg2 ? X16_RX_DATAWIDTH : X20_RX_DATAWIDTH;



//---------- Load Counter ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        load_cnt <= 2'd0;
    else
    
        //---------- Increment Load Counter ----------------
        if ((fsm == FSM_LOAD) && (load_cnt < LOAD_CNT_MAX))
            load_cnt <= load_cnt + 2'd1;
            
        //---------- Hold Load Counter ---------------------
        else if ((fsm == FSM_LOAD) && (load_cnt == LOAD_CNT_MAX))
            load_cnt <= load_cnt;
            
        //---------- Reset Load Counter --------------------
        else
            load_cnt <= 2'd0;
        
end 



//---------- Update DRP Address and Data ---------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        addr_reg <=  9'd0;
        di_reg   <= 16'd0;
        end
    else
        begin
        
        case (index)
        
        //--------------------------------------------------     
        1'd0 :
            begin        
            addr_reg <= ADDR_RX_DATAWIDTH;
            di_reg   <= (do_reg2 & MASK_RX_DATAWIDTH) | data_rx_datawidth;
            end              
            
        //--------------------------------------------------
        default : 
            begin
            addr_reg <=  9'd0;
            di_reg   <= 16'd0;
            end
            
        endcase
        
        end
        
end  



//---------- PIPE DRP FSM ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        fsm   <= FSM_IDLE;
        index <= 5'd0;
        done  <= 1'd0;
        end
    else
        begin
        
        case (fsm)

        //---------- Idle State ----------------------------
        FSM_IDLE :  
          
            begin
            //---------- Reset or Rate Change --------------
            if (start_reg2)
                begin
                fsm   <= FSM_LOAD;
                index <= 5'd0;
                done  <= 1'd0; 
                end
            //---------- Idle ------------------------------
            else       
                begin
                fsm   <= FSM_IDLE;
                index <= 5'd0;
                done  <= 1'd1;
                end 
            end    
            
        //---------- Load DRP Address  ---------------------
        FSM_LOAD :
        
            begin
            fsm   <= (load_cnt == LOAD_CNT_MAX) ? FSM_READ : FSM_LOAD;
            index <= index;

            done  <= 1'd0;
            end  
            
        //---------- Read DRP ------------------------------
        FSM_READ :
        
            begin
            fsm   <= FSM_RRDY;
            index <= index;
            done  <= 1'd0;
            end
            
        //---------- Read DRP Ready ------------------------
        FSM_RRDY :    
        
            begin
            fsm   <= rdy_reg2 ? FSM_WRITE : FSM_RRDY;
            index <= index;
            done  <= 1'd0;
            end
  
            
        //---------- Write DRP -----------------------------
        FSM_WRITE :    
        
            begin
            fsm   <= FSM_WRDY;
            index <= index;
            done  <= 1'd0;
            end       
            
        //---------- Write DRP Ready -----------------------
        FSM_WRDY :    
        
            begin
            fsm   <= rdy_reg2 ? FSM_DONE : FSM_WRDY;
            index <= index;
            done  <= 1'd0;
            end        
             
        //---------- DRP Done ------------------------------
        FSM_DONE :
        
            begin
            if (index == INDEX_MAX)
                begin
                fsm   <= FSM_IDLE;
                index <= 5'd0;
                done  <= 1'd0;
                end
            else       
                begin
                fsm   <= FSM_LOAD;
                index <= index + 5'd1;
                done  <= 1'd0;
                end
            end     
              
        //---------- Default State -------------------------
        default :
        
            begin      
            fsm   <= FSM_IDLE;
            index <= 5'd0;
            done  <= 1'd0;
            end
            
        endcase
        
        end
        
end 



//---------- PIPE DRP Output ---------------------------------------------------
assign DRP_ADDR = addr_reg;
assign DRP_EN   = (fsm == FSM_READ) || (fsm == FSM_WRITE);
assign DRP_DI   = di_reg;
assign DRP_WE   = (fsm == FSM_WRITE);
assign DRP_DONE = done;
assign DRP_FSM  = fsm;



endmodule



`timescale 1ns/1ps
module model_ap2_tst_pipe_drp #
(

    parameter PCIE_GT_DEVICE       = "GTX",                                     // PCIe GT device
    parameter PCIE_USE_MODE        = "3.0",                                     // PCIe use mode
    parameter PCIE_ASYNC_EN        = "FALSE",                                   // PCIe async mode
    parameter PCIE_PLL_SEL         = "CPLL",                                    // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_AUX_CDR_GEN3_EN = "TRUE",                                    // PCIe AUX CDR Gen3 enable
    parameter PCIE_TXBUF_EN        = "FALSE",                                   // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_RXBUF_EN        = "TRUE",                                    // PCIe RX buffer enable for Gen3      only
    parameter PCIE_TXSYNC_MODE     = 0,                                         // PCIe TX sync mode
    parameter PCIE_RXSYNC_MODE     = 0,                                         // PCIe RX sync mode
    parameter LOAD_CNT_MAX         = 2'd1,                                      // Load max count
    parameter INDEX_MAX            = 5'd21                                      // Index max count
    
)

(
    
    //---------- Input -------------------------------------
    input               DRP_CLK,
    input               DRP_RST_N,
    input               DRP_GTXRESET,
    input       [ 1:0]  DRP_RATE,
    input               DRP_X16X20_MODE,
    input               DRP_X16,
    input               DRP_START,
    input       [15:0]  DRP_DO,
    input               DRP_RDY,
    
    //---------- Output ------------------------------------
    output      [ 8:0]  DRP_ADDR,
    output              DRP_EN,  
    output      [15:0]  DRP_DI,   
    output              DRP_WE,
    output              DRP_DONE,
    output      [ 2:0]  DRP_FSM
    
);

    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gtxreset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16x20_mode_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gtxreset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rate_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16x20_mode_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 x16_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg2;
    
    //---------- Internal Signals --------------------------
    reg         [ 1:0]  load_cnt =  2'd0;
    reg         [ 4:0]  index    =  5'd0;
    reg                 mode     =  1'd0;
    reg         [ 8:0]  addr_reg =  9'd0;
    reg         [15:0]  di_reg   = 16'd0;
    
    //---------- Output Registers --------------------------
    reg                 done     =  1'd0;
    reg         [ 2:0]  fsm      =  0;      
                        
    //---------- DRP Address -------------------------------
    //  DRP access for *RXCDR_EIDLE includes 
    //    - [11] RXCDR_HOLD_DURING_EIDLE
    //    - [12] RXCDR_FR_RESET_ON_EIDLE
    //    - [13] RXCDR_PH_RESET_ON_EIDLE
    //------------------------------------------------------
    localparam          ADDR_PCS_RSVD_ATTR        = 9'h06F;
    localparam          ADDR_TXOUT_DIV            = 9'h088;
    localparam          ADDR_RXOUT_DIV            = 9'h088;
    localparam          ADDR_TX_DATA_WIDTH        = 9'h06B;            
    localparam          ADDR_TX_INT_DATAWIDTH     = 9'h06B;         
    localparam          ADDR_RX_DATA_WIDTH        = 9'h011;            
    localparam          ADDR_RX_INT_DATAWIDTH     = 9'h011;              
    localparam          ADDR_TXBUF_EN             = 9'h01C;           
    localparam          ADDR_RXBUF_EN             = 9'h09D;
    localparam          ADDR_TX_XCLK_SEL          = 9'h059;
    localparam          ADDR_RX_XCLK_SEL          = 9'h059;                 
    localparam          ADDR_CLK_CORRECT_USE      = 9'h044; 
    localparam          ADDR_TX_DRIVE_MODE        = 9'h019;
    localparam          ADDR_RXCDR_EIDLE          = 9'h0A7;  
    localparam          ADDR_RX_DFE_LPM_EIDLE     = 9'h01E;
    localparam          ADDR_PMA_RSV_A            = 9'h099;
    localparam          ADDR_PMA_RSV_B            = 9'h09A;
    localparam          ADDR_RXCDR_CFG_A          = 9'h0A8;
    localparam          ADDR_RXCDR_CFG_B          = 9'h0A9;
    localparam          ADDR_RXCDR_CFG_C          = 9'h0AA;
    localparam          ADDR_RXCDR_CFG_D          = 9'h0AB;
    localparam          ADDR_RXCDR_CFG_E          = 9'h0AC;
    localparam          ADDR_RXCDR_CFG_F          = 9'h0AD;  // GTH only
    
    //---------- DRP Mask ----------------------------------
    localparam          MASK_PCS_RSVD_ATTR        = 16'b1111111111111001;  // Unmask bit [ 2: 1]
    localparam          MASK_TXOUT_DIV            = 16'b1111111110001111;  // Unmask bit [ 6: 4]
    localparam          MASK_RXOUT_DIV            = 16'b1111111111111000;  // Unmask bit [ 2: 0]
    localparam          MASK_TX_DATA_WIDTH        = 16'b1111111111111000;  // Unmask bit [ 2: 0]   
    localparam          MASK_TX_INT_DATAWIDTH     = 16'b1111111111101111;  // Unmask bit [    4]
    localparam          MASK_RX_DATA_WIDTH        = 16'b1100011111111111;  // Unmask bit [13:11]  
    localparam          MASK_X16X20_RX_DATA_WIDTH = 16'b1111011111111111;  // Unmask bit [   11] // for x16 or x20 mode only 
    localparam          MASK_RX_INT_DATAWIDTH     = 16'b1011111111111111;  // Unmask bit [   14]  
    localparam          MASK_TXBUF_EN             = 16'b1011111111111111;  // Unmask bit [   14]  
    localparam          MASK_RXBUF_EN             = 16'b1111111111111101;  // Unmask bit [    1] 
    localparam          MASK_TX_XCLK_SEL          = 16'b1111111101111111;  // Unmask bit [    7]    
    localparam          MASK_RX_XCLK_SEL          = 16'b1111111110111111;  // Unmask bit [    6]       
    localparam          MASK_CLK_CORRECT_USE      = 16'b1011111111111111;  // Unmask bit [   14]
    localparam          MASK_TX_DRIVE_MODE        = 16'b1111111111100000;  // Unmask bit [  4:0]      
    localparam          MASK_RXCDR_EIDLE          = 16'b1111011111111111;  // Unmask bit [   11]  
    localparam          MASK_RX_DFE_LPM_EIDLE     = 16'b1011111111111111;  // Unmask bit [   14] 
    localparam          MASK_PMA_RSV_A            = 16'b0000000000000000;  // Unmask bit [15: 0]
    localparam          MASK_PMA_RSV_B            = 16'b0000000000000000;  // Unmask bit [15: 0]
    localparam          MASK_RXCDR_CFG_A          = 16'b0000000000000000;  // Unmask bit [15: 0]
    localparam          MASK_RXCDR_CFG_B          = 16'b0000000000000000;  // Unmask bit [15: 0]
    localparam          MASK_RXCDR_CFG_C          = 16'b0000000000000000;  // Unmask bit [15: 0]    
    localparam          MASK_RXCDR_CFG_D          = 16'b0000000000000000;  // Unmask bit [15: 0]  
    localparam          MASK_RXCDR_CFG_E_GTX      = 16'b1111111100000000;  // Unmask bit [ 7: 0]   
    localparam          MASK_RXCDR_CFG_E_GTH      = 16'b0000000000000000;  // Unmask bit [15: 0] 
    localparam          MASK_RXCDR_CFG_F_GTX      = 16'b1111111111111111;  // Unmask bit [     ] 
    localparam          MASK_RXCDR_CFG_F_GTH      = 16'b1111111111111000;  // Unmask bit [ 2: 0]
         
    //---------- DRP Data for PCIe Gen1 and Gen2 -----------
    localparam          GEN12_TXOUT_DIV           = (PCIE_PLL_SEL == "QPLL") ? 16'b0000000000100000 : 16'b0000000000010000;  // Divide by 4 or 2
    localparam          GEN12_RXOUT_DIV           = (PCIE_PLL_SEL == "QPLL") ? 16'b0000000000000010 : 16'b0000000000000001;  // Divide by 4 or 2
    localparam          GEN12_TX_DATA_WIDTH       = 16'b0000000000000011;  // 2-byte (16-bit) external data width   
    localparam          GEN12_TX_INT_DATAWIDTH    = 16'b0000000000000000;  // 2-byte (20-bit) internal data width
    localparam          GEN12_RX_DATA_WIDTH       = 16'b0001100000000000;  // 2-byte (16-bit) external data width
    localparam          GEN12_RX_INT_DATAWIDTH    = 16'b0000000000000000;  // 2-byte (20-bit) internal data width
    localparam          GEN12_TXBUF_EN            = 16'b0100000000000000;  // Use TX buffer if PCIE_TXBUF_EN == "TRUE"
    localparam          GEN12_RXBUF_EN            = 16'b0000000000000010;  // Use RX buffer 
    localparam          GEN12_TX_XCLK_SEL         = 16'b0000000000000000;  // Use TXOUT if PCIE_TXBUF_EN == "TRUE"
    localparam          GEN12_RX_XCLK_SEL         = 16'b0000000000000000;  // Use RXREC  
    localparam          GEN12_CLK_CORRECT_USE     = 16'b0100000000000000;  // Use clock correction
    localparam          GEN12_TX_DRIVE_MODE       = 16'b0000000000000001;  // Use PIPE   Gen1 and Gen2 mode    
    localparam          GEN12_RXCDR_EIDLE         = 16'b0000100000000000;  // Hold RXCDR during electrical idle 
    localparam          GEN12_RX_DFE_LPM_EIDLE    = 16'b0100000000000000;  // Hold RX DFE or LPM during electrical idle
    localparam          GEN12_PMA_RSV_A_GTX       = 16'b1000010010000000;  // 16'h8480
    localparam          GEN12_PMA_RSV_B_GTX       = 16'b0000000000000001;  // 16'h0001
    localparam          GEN12_PMA_RSV_A_GTH       = 16'b0000000000001000;  // 16'h0008
    localparam          GEN12_PMA_RSV_B_GTH       = 16'b0000000000000000;  // 16'h0000
    //----------
    localparam          GEN12_RXCDR_CFG_A_GTX     = 16'h0020;              // 16'h0020
    localparam          GEN12_RXCDR_CFG_B_GTX     = 16'h1020;              // 16'h1020
    localparam          GEN12_RXCDR_CFG_C_GTX     = 16'h23FF;              // 16'h23FF
    localparam          GEN12_RXCDR_CFG_D_GTX_S   = 16'h0000;              // 16'h0000 Sync
    localparam          GEN12_RXCDR_CFG_D_GTX_A   = 16'h8000;              // 16'h8000 Async    
    localparam          GEN12_RXCDR_CFG_E_GTX     = 16'h0003;              // 16'h0003
    localparam          GEN12_RXCDR_CFG_F_GTX     = 16'h0000;              // 16'h0000
    //----------
    localparam          GEN12_RXCDR_CFG_A_GTH_S   = 16'h0018;              // 16'h0018 Sync
    localparam          GEN12_RXCDR_CFG_A_GTH_A   = 16'h8018;              // 16'h8018 Async
    localparam          GEN12_RXCDR_CFG_B_GTH     = 16'hC208;              // 16'hC208
    localparam          GEN12_RXCDR_CFG_C_GTH     = 16'h2000;              // 16'h2000
    localparam          GEN12_RXCDR_CFG_D_GTH     = 16'h07FE;              // 16'h07FE
    localparam          GEN12_RXCDR_CFG_E_GTH     = 16'h0020;              // 16'h0020
    localparam          GEN12_RXCDR_CFG_F_GTH     = 16'h0000;              // 16'h0000  
    
    //---------- DRP Data for PCIe Gen3 --------------------                 
    localparam          GEN3_TXOUT_DIV            = 16'b0000000000000000;  // Divide by 1
    localparam          GEN3_RXOUT_DIV            = 16'b0000000000000000;  // Divide by 1
    localparam          GEN3_TX_DATA_WIDTH        = 16'b0000000000000100;  // 4-byte (32-bit) external data width                     
    localparam          GEN3_TX_INT_DATAWIDTH     = 16'b0000000000010000;  // 4-byte (32-bit) internal data width               
    localparam          GEN3_RX_DATA_WIDTH        = 16'b0010000000000000;  // 4-byte (32-bit) external data width                  
    localparam          GEN3_RX_INT_DATAWIDTH     = 16'b0100000000000000;  // 4-byte (32-bit) internal data width               
    localparam          GEN3_TXBUF_EN             = 16'b0000000000000000;  // Bypass TX buffer 
    localparam          GEN3_RXBUF_EN             = 16'b0000000000000000;  // Bypass RX buffer  
    localparam          GEN3_TX_XCLK_SEL          = 16'b0000000010000000;  // Use TXUSR  
    localparam          GEN3_RX_XCLK_SEL          = 16'b0000000001000000;  // Use RXUSR                         
    localparam          GEN3_CLK_CORRECT_USE      = 16'b0000000000000000;  // Bypass clock correction  
    localparam          GEN3_TX_DRIVE_MODE        = 16'b0000000000000010;  // Use PIPE Gen3 mode   
    localparam          GEN3_RXCDR_EIDLE          = 16'b0000000000000000;  // Disable Hold RXCDR during electrical idle 
    localparam          GEN3_RX_DFE_LPM_EIDLE     = 16'b0000000000000000;  // Disable RX DFE or LPM during electrical idle   
    localparam          GEN3_PMA_RSV_A_GTX        = 16'b0111000010000000;  // 16'h7080
    localparam          GEN3_PMA_RSV_B_GTX        = 16'b0000000000011110;  // 16'h001E
    localparam          GEN3_PMA_RSV_A_GTH        = 16'b0000000000001000;  // 16'h0008
    localparam          GEN3_PMA_RSV_B_GTH        = 16'b0000000000000000;  // 16'h0000   
    //---------- 
    localparam          GEN3_RXCDR_CFG_A_GTX      = 16'h0080;              // 16'h0080
    localparam          GEN3_RXCDR_CFG_B_GTX      = 16'h1010;              // 16'h1010
    localparam          GEN3_RXCDR_CFG_C_GTX      = 16'h0BFF;              // 16'h0BFF
    localparam          GEN3_RXCDR_CFG_D_GTX_S    = 16'h0000;              // 16'h0000 Sync
    localparam          GEN3_RXCDR_CFG_D_GTX_A    = 16'h8000;              // 16'h8000 Async    
    localparam          GEN3_RXCDR_CFG_E_GTX      = 16'h000B;              // 16'h000B
    localparam          GEN3_RXCDR_CFG_F_GTX      = 16'h0000;              // 16'h0000
    //----------                                 
  //localparam          GEN3_RXCDR_CFG_A_GTH_S    = 16'h0018;              // 16'h0018 Sync
  //localparam          GEN3_RXCDR_CFG_A_GTH_A    = 16'h8018;              // 16'h8018 Async
  //localparam          GEN3_RXCDR_CFG_B_GTH      = 16'hC208;              // 16'hC848
  //localparam          GEN3_RXCDR_CFG_C_GTH      = 16'h2000;              // 16'h1000
  //localparam          GEN3_RXCDR_CFG_D_GTH      = 16'h07FE;              // 16'h07FE v1.0 silicon
  //localparam          GEN3_RXCDR_CFG_D_GTH_AUX  = 16'h0FFE;              // 16'h07FE v2.0 silicon, [62:59] AUX CDR configuration
  //localparam          GEN3_RXCDR_CFG_E_GTH      = 16'h0020;              // 16'h0010
  //localparam          GEN3_RXCDR_CFG_F_GTH      = 16'h0000;              // 16'h0000 v1.0 silicon
  //localparam          GEN3_RXCDR_CFG_F_GTH_AUX  = 16'h0002;              // 16'h0000 v2.0 silicon, [81] AUX CDR enable
    //----------                                 
    localparam          GEN3_RXCDR_CFG_A_GTH_S    = 16'h0018;              // 16'h0018 Sync
    localparam          GEN3_RXCDR_CFG_A_GTH_A    = 16'h8018;              // 16'h8018 Async
    localparam          GEN3_RXCDR_CFG_B_GTH      = 16'hC848;              // 16'hC848
    localparam          GEN3_RXCDR_CFG_C_GTH      = 16'h1000;              // 16'h1000
    localparam          GEN3_RXCDR_CFG_D_GTH      = 16'h07FE;              // 16'h07FE v1.0 silicon
    localparam          GEN3_RXCDR_CFG_D_GTH_AUX  = 16'h0FFE;              // 16'h07FE v2.0 silicon, [62:59] AUX CDR configuration
    localparam          GEN3_RXCDR_CFG_E_GTH      = 16'h0010;              // 16'h0010
    localparam          GEN3_RXCDR_CFG_F_GTH      = 16'h0000;              // 16'h0000 v1.0 silicon
    localparam          GEN3_RXCDR_CFG_F_GTH_AUX  = 16'h0002;              // 16'h0000 v2.0 silicon, [81] AUX CDR enable
      
    //---------- DRP Data for PCIe Gen1, Gen2 and Gen3 -----    
    localparam          GEN123_PCS_RSVD_ATTR_A    = 16'b0000000000000000;  // Auto TX and RX sync mode
    localparam          GEN123_PCS_RSVD_ATTR_M_TX = 16'b0000000000000010;  // Manual TX sync mode
    localparam          GEN123_PCS_RSVD_ATTR_M_RX = 16'b0000000000000100;  // Manual RX sync mode
      
    //---------- DRP Data for x16 --------------------------
    localparam          X16_RX_DATAWIDTH   = 16'b0000000000000000;  // 2-byte (16-bit) internal data width
    
    //---------- DRP Data for x20 --------------------------                                  
    localparam          X20_RX_DATAWIDTH   = 16'b0000100000000000;  // 2-byte (20-bit) internal data width       
      
    //---------- DRP Data ----------------------------------     
    wire        [15:0]  data_txout_div;
    wire        [15:0]  data_rxout_div;
    wire        [15:0]  data_tx_data_width;               
    wire        [15:0]  data_tx_int_datawidth;            
    wire        [15:0]  data_rx_data_width;               
    wire        [15:0]  data_rx_int_datawidth;                
    wire        [15:0]  data_txbuf_en;        
    wire        [15:0]  data_rxbuf_en;        
    wire        [15:0]  data_tx_xclk_sel;
    wire        [15:0]  data_rx_xclk_sel;            
    wire        [15:0]  data_clk_correction_use; 
    wire        [15:0]  data_tx_drive_mode;
    wire        [15:0]  data_rxcdr_eidle;
    wire        [15:0]  data_rx_dfe_lpm_eidle;
    wire        [15:0]  data_pma_rsv_a;
    wire        [15:0]  data_pma_rsv_b;
    
    wire        [15:0]  data_rxcdr_cfg_a;
    wire        [15:0]  data_rxcdr_cfg_b; 
    wire        [15:0]  data_rxcdr_cfg_c;
    wire        [15:0]  data_rxcdr_cfg_d; 
    wire        [15:0]  data_rxcdr_cfg_e;
    wire        [15:0]  data_rxcdr_cfg_f;
        
    wire        [15:0]  data_pcs_rsvd_attr_a;  
    wire        [15:0]  data_pcs_rsvd_attr_m_tx; 
    wire        [15:0]  data_pcs_rsvd_attr_m_rx; 
    wire        [15:0]  data_pcs_rsvd_attr_m;   
                
    wire        [15:0]  data_x16x20_rx_datawidth;    
           
    //---------- FSM ---------------------------------------  
    localparam          FSM_IDLE  = 0;  
    localparam          FSM_LOAD  = 1;                           
    localparam          FSM_READ  = 2;
    localparam          FSM_RRDY  = 3;
    localparam          FSM_WRITE = 4;
    localparam          FSM_WRDY  = 5;    
    localparam          FSM_DONE  = 6;   

    
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        //---------- 1st Stage FF --------------------------
        gtxreset_reg1    <=  1'd0;
        rate_reg1        <=  2'd0;
        x16x20_mode_reg1 <=  1'd0;
        x16_reg1         <=  1'd0;
        do_reg1          <= 16'd0;
        rdy_reg1         <=  1'd0;
        start_reg1       <=  1'd0;
        //---------- 2nd Stage FF --------------------------
        gtxreset_reg2    <=  1'd0;
        rate_reg2        <=  2'd0;
        x16x20_mode_reg2 <=  1'd0;
        x16_reg2         <=  1'd0;
        do_reg2          <= 16'd0;
        rdy_reg2         <=  1'd0;
        start_reg2       <=  1'd0;
        end
        
    else
        begin
        //---------- 1st Stage FF --------------------------
        gtxreset_reg1    <= DRP_GTXRESET;
        rate_reg1        <= DRP_RATE;
        x16x20_mode_reg1 <= DRP_X16X20_MODE;
        x16_reg1         <= DRP_X16;
        do_reg1          <= DRP_DO;
        rdy_reg1         <= DRP_RDY;
        start_reg1       <= DRP_START;
        //---------- 2nd Stage FF --------------------------
        gtxreset_reg2    <= gtxreset_reg1;
        rate_reg2        <= rate_reg1;
        x16x20_mode_reg2 <= x16x20_mode_reg1;
        x16_reg2         <= x16_reg1;
        do_reg2          <= do_reg1;
        rdy_reg2         <= rdy_reg1;
        start_reg2       <= start_reg1;
        end
    
end  



//---------- Select DRP Data ---------------------------------------------------
assign data_txout_div          =  (rate_reg2 == 2'd2)                                ? GEN3_TXOUT_DIV        : GEN12_TXOUT_DIV;
assign data_rxout_div          =  (rate_reg2 == 2'd2)                                ? GEN3_RXOUT_DIV        : GEN12_RXOUT_DIV;
assign data_tx_data_width      =  (rate_reg2 == 2'd2)                                ? GEN3_TX_DATA_WIDTH    : GEN12_TX_DATA_WIDTH;
assign data_tx_int_datawidth   =  (rate_reg2 == 2'd2)                                ? GEN3_TX_INT_DATAWIDTH : GEN12_TX_INT_DATAWIDTH;
assign data_rx_data_width      =  (rate_reg2 == 2'd2)                                ? GEN3_RX_DATA_WIDTH    : GEN12_RX_DATA_WIDTH;

assign data_rx_int_datawidth   =  (rate_reg2 == 2'd2)                                ? GEN3_RX_INT_DATAWIDTH : GEN12_RX_INT_DATAWIDTH;

assign data_txbuf_en           = ((rate_reg2 == 2'd2) || (PCIE_TXBUF_EN == "FALSE")) ? GEN3_TXBUF_EN         : GEN12_TXBUF_EN;
assign data_rxbuf_en           = ((rate_reg2 == 2'd2) && (PCIE_RXBUF_EN == "FALSE")) ? GEN3_RXBUF_EN         : GEN12_RXBUF_EN;
assign data_tx_xclk_sel        = ((rate_reg2 == 2'd2) || (PCIE_TXBUF_EN == "FALSE")) ? GEN3_TX_XCLK_SEL      : GEN12_TX_XCLK_SEL;
assign data_rx_xclk_sel        = ((rate_reg2 == 2'd2) && (PCIE_RXBUF_EN == "FALSE")) ? GEN3_RX_XCLK_SEL      : GEN12_RX_XCLK_SEL;
assign data_clk_correction_use =  (rate_reg2 == 2'd2)                                ? GEN3_CLK_CORRECT_USE  : GEN12_CLK_CORRECT_USE;
assign data_tx_drive_mode      =  (rate_reg2 == 2'd2)                                ? GEN3_TX_DRIVE_MODE    : GEN12_TX_DRIVE_MODE;   
assign data_rxcdr_eidle        =  (rate_reg2 == 2'd2)                                ? GEN3_RXCDR_EIDLE      : GEN12_RXCDR_EIDLE;
assign data_rx_dfe_lpm_eidle   =  (rate_reg2 == 2'd2)                                ? GEN3_RX_DFE_LPM_EIDLE : GEN12_RX_DFE_LPM_EIDLE;
assign data_pma_rsv_a          =  (rate_reg2 == 2'd2)                                ? ((PCIE_GT_DEVICE == "GTH") ? GEN3_PMA_RSV_A_GTH  : GEN3_PMA_RSV_A_GTX) :
                                                                                       ((PCIE_GT_DEVICE == "GTH") ? GEN12_PMA_RSV_A_GTH : GEN12_PMA_RSV_A_GTX);
assign data_pma_rsv_b          =  (rate_reg2 == 2'd2)                                ? ((PCIE_GT_DEVICE == "GTH") ? GEN3_PMA_RSV_B_GTH  : GEN3_PMA_RSV_B_GTX) :
                                                                                       ((PCIE_GT_DEVICE == "GTH") ? GEN12_PMA_RSV_B_GTH : GEN12_PMA_RSV_B_GTX);

assign data_rxcdr_cfg_a = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ? ((PCIE_ASYNC_EN == "TRUE") ? GEN3_RXCDR_CFG_A_GTH_A  : GEN3_RXCDR_CFG_A_GTH_S)  : GEN3_RXCDR_CFG_A_GTX) :
                                                ((PCIE_GT_DEVICE == "GTH") ? ((PCIE_ASYNC_EN == "TRUE") ? GEN12_RXCDR_CFG_A_GTH_A : GEN12_RXCDR_CFG_A_GTH_S) : GEN12_RXCDR_CFG_A_GTX);

assign data_rxcdr_cfg_b = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ?  GEN3_RXCDR_CFG_B_GTH  : GEN3_RXCDR_CFG_B_GTX) :
                                                ((PCIE_GT_DEVICE == "GTH") ?  GEN12_RXCDR_CFG_B_GTH : GEN12_RXCDR_CFG_B_GTX);

assign data_rxcdr_cfg_c = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ?  GEN3_RXCDR_CFG_C_GTH  : GEN3_RXCDR_CFG_C_GTX) :
                                                ((PCIE_GT_DEVICE == "GTH") ?  GEN12_RXCDR_CFG_C_GTH : GEN12_RXCDR_CFG_C_GTX);
                                                
assign data_rxcdr_cfg_d = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ?  ((PCIE_AUX_CDR_GEN3_EN == "TRUE") ? GEN3_RXCDR_CFG_D_GTH_AUX : GEN3_RXCDR_CFG_D_GTH) : ((PCIE_ASYNC_EN == "TRUE") ? GEN3_RXCDR_CFG_D_GTX_A : GEN3_RXCDR_CFG_D_GTX_S)) :
                                                ((PCIE_GT_DEVICE == "GTH") ?  GEN12_RXCDR_CFG_D_GTH : ((PCIE_ASYNC_EN == "TRUE") ? GEN3_RXCDR_CFG_D_GTX_A : GEN3_RXCDR_CFG_D_GTX_S));

assign data_rxcdr_cfg_e = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ?  GEN3_RXCDR_CFG_E_GTH  : GEN3_RXCDR_CFG_E_GTX) :
                                                ((PCIE_GT_DEVICE == "GTH") ?  GEN12_RXCDR_CFG_E_GTH : GEN12_RXCDR_CFG_E_GTX);
                                                
assign data_rxcdr_cfg_f = (rate_reg2 == 2'd2) ? ((PCIE_GT_DEVICE == "GTH") ?  ((PCIE_AUX_CDR_GEN3_EN == "TRUE") ? GEN3_RXCDR_CFG_F_GTH_AUX : GEN3_RXCDR_CFG_F_GTH) : GEN3_RXCDR_CFG_F_GTX) :
                                                ((PCIE_GT_DEVICE == "GTH") ?  GEN12_RXCDR_CFG_F_GTH : GEN12_RXCDR_CFG_F_GTX);

assign data_pcs_rsvd_attr_a    = GEN123_PCS_RSVD_ATTR_A;
assign data_pcs_rsvd_attr_m_tx = PCIE_TXSYNC_MODE ? GEN123_PCS_RSVD_ATTR_A : GEN123_PCS_RSVD_ATTR_M_TX;
assign data_pcs_rsvd_attr_m_rx = PCIE_RXSYNC_MODE ? GEN123_PCS_RSVD_ATTR_A : GEN123_PCS_RSVD_ATTR_M_RX;
assign data_pcs_rsvd_attr_m    = data_pcs_rsvd_attr_m_tx | data_pcs_rsvd_attr_m_rx;

assign data_x16x20_rx_datawidth = x16_reg2 ? X16_RX_DATAWIDTH : X20_RX_DATAWIDTH;


//---------- Load Counter ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        load_cnt <= 2'd0;
    else
    
        //---------- Increment Load Counter ----------------
        if ((fsm == FSM_LOAD) && (load_cnt < LOAD_CNT_MAX))
            load_cnt <= load_cnt + 2'd1;
            
        //---------- Hold Load Counter ---------------------
        else if ((fsm == FSM_LOAD) && (load_cnt == LOAD_CNT_MAX))
            load_cnt <= load_cnt;
            
        //---------- Reset Load Counter --------------------
        else
            load_cnt <= 2'd0;
        
end 



//---------- Update DRP Address and Data ---------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        addr_reg <=  9'd0;
        di_reg   <= 16'd0;
        end
    else
        begin
        
        case (index)
        
        //--------------------------------------------------      
        5'd0:     
            begin
            addr_reg <= mode             ? ADDR_PCS_RSVD_ATTR : 
                        x16x20_mode_reg2 ? ADDR_RX_DATA_WIDTH : ADDR_TXOUT_DIV; 
            di_reg   <= mode             ? ((do_reg2 & MASK_PCS_RSVD_ATTR)        | data_pcs_rsvd_attr_a) : 
                        x16x20_mode_reg2 ? ((do_reg2 & MASK_X16X20_RX_DATA_WIDTH) | data_x16x20_rx_datawidth) : 
                                           ((do_reg2 & MASK_TXOUT_DIV)            | data_txout_div);
            end 
            
        //--------------------------------------------------      
        5'd1:    
            begin
            addr_reg <= mode ? ADDR_PCS_RSVD_ATTR : ADDR_RXOUT_DIV;
            di_reg   <= mode ? ((do_reg2 & MASK_PCS_RSVD_ATTR)  | data_pcs_rsvd_attr_m) : 
                               ((do_reg2 & MASK_RXOUT_DIV)      | data_rxout_div);
            end 
            
        //--------------------------------------------------
        5'd2 :
            begin        
            addr_reg <= ADDR_TX_DATA_WIDTH;
            di_reg   <= (do_reg2 & MASK_TX_DATA_WIDTH) | data_tx_data_width;
            end
           
        //--------------------------------------------------    
        5'd3 :
            begin        
            addr_reg <= ADDR_TX_INT_DATAWIDTH;
            di_reg   <= (do_reg2 & MASK_TX_INT_DATAWIDTH) | data_tx_int_datawidth;
            end    
        
        //--------------------------------------------------     
        5'd4 :
            begin
            addr_reg <= ADDR_RX_DATA_WIDTH;
            di_reg   <= (do_reg2 & MASK_RX_DATA_WIDTH) | data_rx_data_width;
            end   
        
        //--------------------------------------------------     
        5'd5 :
            begin        
            addr_reg <= ADDR_RX_INT_DATAWIDTH;
            di_reg   <= (do_reg2 & MASK_RX_INT_DATAWIDTH) | data_rx_int_datawidth;
            end  
  
        //--------------------------------------------------         
        5'd6 :
            begin        
            addr_reg <= ADDR_TXBUF_EN;
            di_reg   <= (do_reg2 & MASK_TXBUF_EN) | data_txbuf_en;
            end   
        
        //--------------------------------------------------         
        5'd7 :
            begin        
            addr_reg <= ADDR_RXBUF_EN;
            di_reg   <= (do_reg2 & MASK_RXBUF_EN) | data_rxbuf_en;
            end   
        
        //--------------------------------------------------         
        5'd8 :
            begin        
            addr_reg <= ADDR_TX_XCLK_SEL;
            di_reg   <= (do_reg2 & MASK_TX_XCLK_SEL) | data_tx_xclk_sel;
            end   
        
        //--------------------------------------------------         
        5'd9 :
            begin        
            addr_reg <= ADDR_RX_XCLK_SEL;
            di_reg   <= (do_reg2 & MASK_RX_XCLK_SEL) | data_rx_xclk_sel;
            end   
        
        //--------------------------------------------------      
        5'd10 :
            begin
            addr_reg <= ADDR_CLK_CORRECT_USE;
            di_reg   <= (do_reg2 & MASK_CLK_CORRECT_USE) | data_clk_correction_use;
            end 

        //--------------------------------------------------      
        5'd11 :
            begin
            addr_reg <= ADDR_TX_DRIVE_MODE;
            di_reg   <= (do_reg2 & MASK_TX_DRIVE_MODE) | data_tx_drive_mode;
            end 
            
        //--------------------------------------------------      
        5'd12 :
            begin
            addr_reg <= ADDR_RXCDR_EIDLE;
            di_reg   <= (do_reg2 & MASK_RXCDR_EIDLE) | data_rxcdr_eidle;
            end 
            
        //--------------------------------------------------      
        5'd13 :
            begin
            addr_reg <= ADDR_RX_DFE_LPM_EIDLE;
            di_reg   <= (do_reg2 & MASK_RX_DFE_LPM_EIDLE) | data_rx_dfe_lpm_eidle;
            end     
            
        //--------------------------------------------------      
        5'd14 :
            begin
            addr_reg <= ADDR_PMA_RSV_A;
            di_reg   <= (do_reg2 & MASK_PMA_RSV_A) | data_pma_rsv_a;
            end  
            
        //--------------------------------------------------      
        5'd15 :
            begin
            addr_reg <= ADDR_PMA_RSV_B;
            di_reg   <= (do_reg2 & MASK_PMA_RSV_B) | data_pma_rsv_b;
            end 

        //--------------------------------------------------      
        5'd16 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_A;
            di_reg   <= (do_reg2 & MASK_RXCDR_CFG_A) | data_rxcdr_cfg_a;
            end 
            
        //--------------------------------------------------      
        5'd17 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_B;
            di_reg   <= (do_reg2 & MASK_RXCDR_CFG_B) | data_rxcdr_cfg_b;
            end 
            
        //--------------------------------------------------      
        5'd18 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_C;
            di_reg   <= (do_reg2 & MASK_RXCDR_CFG_C) | data_rxcdr_cfg_c;
            end                         

        //--------------------------------------------------      
        5'd19 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_D;
            di_reg   <= (do_reg2 & MASK_RXCDR_CFG_D) | data_rxcdr_cfg_d;
            end    
            
        //--------------------------------------------------      
        5'd20 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_E;
            di_reg   <= (do_reg2 & ((PCIE_GT_DEVICE == "GTH") ? MASK_RXCDR_CFG_E_GTH : MASK_RXCDR_CFG_E_GTX)) | data_rxcdr_cfg_e;
            end             
            
        //--------------------------------------------------      
        5'd21 :
            begin
            addr_reg <= ADDR_RXCDR_CFG_F;
            di_reg   <= (do_reg2 & ((PCIE_GT_DEVICE == "GTH") ? MASK_RXCDR_CFG_F_GTH : MASK_RXCDR_CFG_F_GTX)) | data_rxcdr_cfg_f;
            end             
            
        //--------------------------------------------------
        default : 
            begin
            addr_reg <=  9'd0;
            di_reg   <= 16'd0;
            end
            
        endcase
        
        end
        
end  



//---------- PIPE DRP FSM ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        fsm   <= FSM_IDLE;
        index <= 5'd0;
        mode  <= 1'd0;
        done  <= 1'd0;
        end
    else
        begin
        
        case (fsm)

        //---------- Idle State ----------------------------
        FSM_IDLE :  
          
            begin
            //---------- Reset or Rate Change --------------
            if (start_reg2)
                begin
                fsm   <= FSM_LOAD;
                index <= 5'd0;
                mode  <= 1'd0;
                done  <= 1'd0; 
                end
            //---------- GTXRESET --------------------------    
            else if ((gtxreset_reg2 && !gtxreset_reg1) && ((PCIE_TXSYNC_MODE == 0) || (PCIE_RXSYNC_MODE == 0)) && (PCIE_USE_MODE == "1.0"))
                begin
                fsm   <= FSM_LOAD;
                index <= 5'd0;
                mode  <= 1'd1;
                done  <= 1'd0;
                end
            //---------- Idle ------------------------------
            else       
                begin
                fsm   <= FSM_IDLE;
                index <= 5'd0;
                mode  <= 1'd0;
                done  <= 1'd1;
                end 
            end    
            
        //---------- Load DRP Address  ---------------------
        FSM_LOAD :
        
            begin
            fsm   <= (load_cnt == LOAD_CNT_MAX) ? FSM_READ : FSM_LOAD;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end  
            
        //---------- Read DRP ------------------------------
        FSM_READ :
        
            begin
            fsm   <= FSM_RRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end
            
        //---------- Read DRP Ready ------------------------
        FSM_RRDY :    
        
            begin
            fsm   <= rdy_reg2 ? FSM_WRITE : FSM_RRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end
  
            
        //---------- Write DRP -----------------------------
        FSM_WRITE :    
        
            begin
            fsm   <= FSM_WRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end       
            
        //---------- Write DRP Ready -----------------------
        FSM_WRDY :    
        
            begin
            fsm   <= rdy_reg2 ? FSM_DONE : FSM_WRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end        
             
        //---------- DRP Done ------------------------------
        FSM_DONE :
        
            begin
            if ((index == INDEX_MAX) || (mode && (index == 5'd1)) || (x16x20_mode_reg2 && (index == 5'd0)))
                begin
                fsm   <= FSM_IDLE;
                index <= 5'd0;
                mode  <= 1'd0;
                done  <= 1'd0;
                end
            else       
                begin
                fsm   <= FSM_LOAD;
                index <= index + 5'd1;
                mode  <= mode;
                done  <= 1'd0;
                end
            end     
              
        //---------- Default State -------------------------
        default :
        
            begin      
            fsm   <= FSM_IDLE;
            index <= 5'd0;
            mode  <= 1'd0;
            done  <= 1'd0;
            end
            
        endcase
        
        end
        
end 



//---------- PIPE DRP Output ---------------------------------------------------
assign DRP_ADDR = addr_reg;
assign DRP_EN   = (fsm == FSM_READ) || (fsm == FSM_WRITE);
assign DRP_DI   = di_reg;
assign DRP_WE   = (fsm == FSM_WRITE);
assign DRP_DONE = done;
assign DRP_FSM  = fsm;



endmodule




`timescale 1ns/1ps
module model_ap2_tst_pipe_eq #
(
    parameter PCIE_SIM_MODE       = "FALSE",
    parameter PCIE_GT_DEVICE      = "GTX",
    parameter PCIE_RXEQ_MODE_GEN3 = 1
)

(

    //---------- Input -------------------------------------
    input               EQ_CLK,                            
    input               EQ_RST_N,
    input               EQ_GEN3,

    input       [ 1:0]  EQ_TXEQ_CONTROL,    
    input       [ 3:0]  EQ_TXEQ_PRESET,
    input       [ 3:0]  EQ_TXEQ_PRESET_DEFAULT,
    input       [ 5:0]  EQ_TXEQ_DEEMPH_IN,
                                
    input       [ 1:0]  EQ_RXEQ_CONTROL,  
    input       [ 2:0]  EQ_RXEQ_PRESET,
    input       [ 5:0]  EQ_RXEQ_LFFS,  
    input       [ 3:0]  EQ_RXEQ_TXPRESET,
    input               EQ_RXEQ_USER_EN,
    input       [17:0]  EQ_RXEQ_USER_TXCOEFF,
    input               EQ_RXEQ_USER_MODE, 
    
    
    //---------- Output ------------------------------------
    output              EQ_TXEQ_DEEMPH,
    output      [ 4:0]  EQ_TXEQ_PRECURSOR,
    output      [ 6:0]  EQ_TXEQ_MAINCURSOR,
    output      [ 4:0]  EQ_TXEQ_POSTCURSOR,
    output      [17:0]  EQ_TXEQ_DEEMPH_OUT,
    output              EQ_TXEQ_DONE,
    output      [ 5:0]  EQ_TXEQ_FSM,
    
    output      [17:0]  EQ_RXEQ_NEW_TXCOEFF,
    output              EQ_RXEQ_LFFS_SEL,
    output              EQ_RXEQ_ADAPT_DONE,
    output              EQ_RXEQ_DONE, 
    output      [ 5:0]  EQ_RXEQ_FSM

);          

    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg2;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  txeq_control_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 3:0]  txeq_preset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  txeq_deemph_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  txeq_control_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg	      [ 3:0]  txeq_preset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  txeq_deemph_reg2;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rxeq_control_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg	      [ 2:0]  rxeq_preset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  rxeq_lffs_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 3:0]  rxeq_txpreset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_user_en_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [17:0]  rxeq_user_txcoeff_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_user_mode_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 1:0]  rxeq_control_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg	      [ 2:0]  rxeq_preset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  rxeq_lffs_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 3:0]  rxeq_txpreset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_user_en_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [17:0]  rxeq_user_txcoeff_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rxeq_user_mode_reg2;
    
    //---------- Internal Signals --------------------------
    reg         [18:0]  txeq_preset          = 19'd0;          
    reg                 txeq_preset_done     =  1'd0;
    reg         [ 1:0]  txeq_txcoeff_cnt     =  2'd0;
    
    reg         [ 2:0]  rxeq_preset          =  3'd0;
    reg                 rxeq_preset_valid    =  1'd0;
    reg         [ 3:0]  rxeq_txpreset        =  4'd0;
    reg         [17:0]  rxeq_txcoeff         = 18'd0; 
    reg         [ 2:0]  rxeq_cnt             =  3'd0;
    reg         [ 5:0]  rxeq_fs              =  6'd0;
    reg         [ 5:0]  rxeq_lf              =  6'd0;
    reg                 rxeq_new_txcoeff_req =  1'd0;
   
    //---------- Output Registers --------------------------     
    reg         [18:0]  txeq_txcoeff        = 19'd0;
    reg                 txeq_done           =  1'd0;
    reg         [ 5:0]  fsm_tx              =  6'd0;
   
    reg         [17:0]  rxeq_new_txcoeff    = 18'd0;
    reg                 rxeq_lffs_sel       =  1'd0;
    reg                 rxeq_adapt_done_reg =  1'd0;
    reg                 rxeq_adapt_done     =  1'd0;
    reg                 rxeq_done           =  1'd0; 
    reg         [ 5:0]  fsm_rx              =  6'd0;    
    
    //---------- RXEQ Eye Scan Module Output ---------------
    wire                rxeqscan_lffs_sel;
    wire                rxeqscan_preset_done;
    wire        [17:0]  rxeqscan_new_txcoeff;
    wire                rxeqscan_new_txcoeff_done;
    wire                rxeqscan_adapt_done;
                  
    //---------- FSM ---------------------------------------   
    localparam          FSM_TXEQ_IDLE            = 6'b000001; 
    localparam          FSM_TXEQ_PRESET          = 6'b000010;                                     
    localparam          FSM_TXEQ_TXCOEFF         = 6'b000100;
    localparam          FSM_TXEQ_REMAP           = 6'b001000;
    localparam          FSM_TXEQ_QUERY           = 6'b010000;                                     
    localparam          FSM_TXEQ_DONE            = 6'b100000;
                                          
    localparam          FSM_RXEQ_IDLE            = 6'b000001; 
    localparam          FSM_RXEQ_PRESET          = 6'b000010;                                     
    localparam          FSM_RXEQ_TXCOEFF         = 6'b000100;
    localparam          FSM_RXEQ_LF              = 6'b001000;
    localparam          FSM_RXEQ_NEW_TXCOEFF_REQ = 6'b010000;                                  
    localparam          FSM_RXEQ_DONE            = 6'b100000;
                
    //---------- TXEQ Presets Look-up Table ----------------
    // TXPRECURSOR  = Coefficient range between  0 and 20 units 
    // TXMAINCURSOR = Coefficient range between 29 and 80 units
    // TXPOSTCURSOR = Coefficient range between  0 and 31 units
    //------------------------------------------------------
    // Actual    Full Swing    (FS) = 80
    // Actual    Low Frequency (LF) = 29
    // Advertise Full Swing    (FS) = 40
    // Advertise Low Frequency (LF) = 15
    //------------------------------------------------------
    // Pre-emphasis  = 20 log [80 - (2 * TXPRECURSOR)] / 80], assuming no de-emphasis
    // Main-emphasis = 80 - (TXPRECURSOR + TXPOSTCURSOR)
    // De-emphasis   = 20 log [80 - (2 *  TXPOSTCURSOR)] / 80], assuming no pre-emphasis
    //------------------------------------------------------    
    // Note:  TXMAINCURSOR calculated internally in GT
    //------------------------------------------------------                           
    localparam          TXPRECURSOR_00  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_00 = 7'd60;                                
    localparam          TXPOSTCURSOR_00 = 6'd20;            // -6.0 +/- 1 dB
    
    localparam          TXPRECURSOR_01  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_01 = 7'd68;            // added 1 to compensate decimal                                
    localparam          TXPOSTCURSOR_01 = 6'd13;            // -3.5 +/- 1 dB
    
    localparam          TXPRECURSOR_02  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_02 = 7'd64;                                
    localparam          TXPOSTCURSOR_02 = 6'd16;            // -4.4 +/- 1.5 dB
    
    localparam          TXPRECURSOR_03  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_03 = 7'd70;                                
    localparam          TXPOSTCURSOR_03 = 6'd10;            // -2.5 +/- 1 dB

    localparam          TXPRECURSOR_04  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_04 = 7'd80;                                
    localparam          TXPOSTCURSOR_04 = 6'd0;             //  0.0 dB
    
    localparam          TXPRECURSOR_05  = 6'd8;             // -1.9 +/- 1 dB
    localparam          TXMAINCURSOR_05 = 7'd72;                                
    localparam          TXPOSTCURSOR_05 = 6'd0;             //  0.0 dB
    
    localparam          TXPRECURSOR_06  = 6'd10;            // -2.5 +/- 1 dB
    localparam          TXMAINCURSOR_06 = 7'd70;                                
    localparam          TXPOSTCURSOR_06 = 6'd0;             //  0.0 dB
    
    localparam          TXPRECURSOR_07  = 6'd8;             // -3.5 +/- 1 dB
    localparam          TXMAINCURSOR_07 = 7'd56;                                
    localparam          TXPOSTCURSOR_07 = 6'd16;            // -6.0 +/- 1 dB
        
    localparam          TXPRECURSOR_08  = 6'd10;            // -3.5 +/- 1 dB
    localparam          TXMAINCURSOR_08 = 7'd60;                                
    localparam          TXPOSTCURSOR_08 = 6'd10;            // -3.5 +/- 1 dB
    
    localparam          TXPRECURSOR_09  = 6'd13;            // -3.5 +/- 1 dB
    localparam          TXMAINCURSOR_09 = 7'd68;            //  added 1 to compensate decimal                  
    localparam          TXPOSTCURSOR_09 = 6'd0;             //  0.0 dB
    
    localparam          TXPRECURSOR_10  = 6'd0;             //  0.0 dB
    localparam          TXMAINCURSOR_10 = 7'd56;            //  added 1 to compensate decimal                     
    localparam          TXPOSTCURSOR_10 = 6'd25;            //  9.5 +/- 1 dB, updated for coefficient rules
    
    
    
//---------- Input FF ----------------------------------------------------------
always @ (posedge EQ_CLK)
begin

    if (!EQ_RST_N)
        begin   
        //---------- 1st Stage FF --------------------------  
        gen3_reg1              <=  1'd0;
                                  
        txeq_control_reg1      <=  2'd0;
        txeq_preset_reg1       <=  4'd0;
        txeq_deemph_reg1       <=  6'd1;
                                  
        rxeq_control_reg1      <=  2'd0;
        rxeq_preset_reg1       <=  3'd0;
        rxeq_lffs_reg1         <=  6'd0;
        rxeq_txpreset_reg1     <=  4'd0;
        rxeq_user_en_reg1      <=  1'd0;
        rxeq_user_txcoeff_reg1 <= 18'd0;
        rxeq_user_mode_reg1    <=  1'd0;
        //---------- 2nd Stage FF --------------------------
        gen3_reg2              <=  1'd0;
                                   
        txeq_control_reg2      <=  2'd0;
        txeq_preset_reg2       <=  4'd0;
        txeq_deemph_reg2       <=  6'd1;
                                   
        rxeq_control_reg2      <=  2'd0;
        rxeq_preset_reg2       <=  3'd0;
        rxeq_lffs_reg2         <=  6'd0;
        rxeq_txpreset_reg2     <=  4'd0;
        rxeq_user_en_reg2      <=  1'd0;
        rxeq_user_txcoeff_reg2 <= 18'd0;
        rxeq_user_mode_reg2    <=  1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF -------------------------- 
        gen3_reg1              <= EQ_GEN3;
                               
        txeq_control_reg1      <= EQ_TXEQ_CONTROL;
        txeq_preset_reg1       <= EQ_TXEQ_PRESET;
        txeq_deemph_reg1       <= EQ_TXEQ_DEEMPH_IN;
                               
        rxeq_control_reg1      <= EQ_RXEQ_CONTROL;
        rxeq_preset_reg1       <= EQ_RXEQ_PRESET;
        rxeq_lffs_reg1         <= EQ_RXEQ_LFFS;
        rxeq_txpreset_reg1     <= EQ_RXEQ_TXPRESET;
        rxeq_user_en_reg1      <= EQ_RXEQ_USER_EN;
        rxeq_user_txcoeff_reg1 <= EQ_RXEQ_USER_TXCOEFF;
        rxeq_user_mode_reg1    <= EQ_RXEQ_USER_MODE;
        //---------- 2nd Stage FF -------------------------- 
        gen3_reg2              <= gen3_reg1;
                               
        txeq_control_reg2      <= txeq_control_reg1;
        txeq_preset_reg2       <= txeq_preset_reg1;
        txeq_deemph_reg2       <= txeq_deemph_reg1;
                               
        rxeq_control_reg2      <= rxeq_control_reg1;
        rxeq_preset_reg2       <= rxeq_preset_reg1;
        rxeq_lffs_reg2         <= rxeq_lffs_reg1;
        rxeq_txpreset_reg2     <= rxeq_txpreset_reg1;
        rxeq_user_en_reg2      <= rxeq_user_en_reg1;
        rxeq_user_txcoeff_reg2 <= rxeq_user_txcoeff_reg1;
        rxeq_user_mode_reg2    <= rxeq_user_mode_reg1;
        end
        
end       



//---------- TXEQ Preset -------------------------------------------------------
always @ (posedge EQ_CLK)
begin

    if (!EQ_RST_N)
        begin
        
        //---------- Select TXEQ Preset ----------------
        case (EQ_TXEQ_PRESET_DEFAULT)
        4'd0    : txeq_preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};
        4'd1    : txeq_preset <= {TXPOSTCURSOR_01, TXMAINCURSOR_01, TXPRECURSOR_01};
        4'd2    : txeq_preset <= {TXPOSTCURSOR_02, TXMAINCURSOR_02, TXPRECURSOR_02};
        4'd3    : txeq_preset <= {TXPOSTCURSOR_03, TXMAINCURSOR_03, TXPRECURSOR_03};
        4'd4    : txeq_preset <= {TXPOSTCURSOR_04, TXMAINCURSOR_04, TXPRECURSOR_04};
        4'd5    : txeq_preset <= {TXPOSTCURSOR_05, TXMAINCURSOR_05, TXPRECURSOR_05};
        4'd6    : txeq_preset <= {TXPOSTCURSOR_06, TXMAINCURSOR_06, TXPRECURSOR_06};
        4'd7    : txeq_preset <= {TXPOSTCURSOR_07, TXMAINCURSOR_07, TXPRECURSOR_07};
        4'd8    : txeq_preset <= {TXPOSTCURSOR_08, TXMAINCURSOR_08, TXPRECURSOR_08};      
        4'd9    : txeq_preset <= {TXPOSTCURSOR_09, TXMAINCURSOR_09, TXPRECURSOR_09};   
        4'd10   : txeq_preset <= {TXPOSTCURSOR_10, TXMAINCURSOR_10, TXPRECURSOR_10};                 
        default : txeq_preset <= 19'd4;     
        endcase
        	   
        txeq_preset_done <=  1'd0;
        end                    
    else
        begin   
        if (fsm_tx == FSM_TXEQ_PRESET)
            begin
            
            //---------- Select TXEQ Preset ----------------
            case (txeq_preset_reg2)
            4'd0    : txeq_preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};
            4'd1    : txeq_preset <= {TXPOSTCURSOR_01, TXMAINCURSOR_01, TXPRECURSOR_01};
            4'd2    : txeq_preset <= {TXPOSTCURSOR_02, TXMAINCURSOR_02, TXPRECURSOR_02};
            4'd3    : txeq_preset <= {TXPOSTCURSOR_03, TXMAINCURSOR_03, TXPRECURSOR_03};
            4'd4    : txeq_preset <= {TXPOSTCURSOR_04, TXMAINCURSOR_04, TXPRECURSOR_04};
            4'd5    : txeq_preset <= {TXPOSTCURSOR_05, TXMAINCURSOR_05, TXPRECURSOR_05};
            4'd6    : txeq_preset <= {TXPOSTCURSOR_06, TXMAINCURSOR_06, TXPRECURSOR_06};
            4'd7    : txeq_preset <= {TXPOSTCURSOR_07, TXMAINCURSOR_07, TXPRECURSOR_07};
            4'd8    : txeq_preset <= {TXPOSTCURSOR_08, TXMAINCURSOR_08, TXPRECURSOR_08};      
            4'd9    : txeq_preset <= {TXPOSTCURSOR_09, TXMAINCURSOR_09, TXPRECURSOR_09}; 
            4'd10   : txeq_preset <= {TXPOSTCURSOR_10, TXMAINCURSOR_10, TXPRECURSOR_10};                   
            default : txeq_preset <= 19'd4;     
        	   endcase
        
            txeq_preset_done <= 1'd1;
            end
        else
            begin
            txeq_preset      <= txeq_preset;
            txeq_preset_done <= 1'd0;
            end
        end
        
end     



//---------- TXEQ FSM ----------------------------------------------------------
always @ (posedge EQ_CLK)
begin

    if (!EQ_RST_N)
        begin
        fsm_tx           <=  FSM_TXEQ_IDLE; 
        txeq_txcoeff     <= 19'd0;
        txeq_txcoeff_cnt <=  2'd0;
        txeq_done        <=  1'd0;
        end                    
    else
        begin
        
        case (fsm_tx)
        
        //---------- Idle State ----------------------------
        FSM_TXEQ_IDLE :
        
            begin
            
            case (txeq_control_reg2)
            
            //---------- Idle ------------------------------
            2'd0    :
                begin
                fsm_tx           <= FSM_TXEQ_IDLE; 
                txeq_txcoeff     <= txeq_txcoeff;
                txeq_txcoeff_cnt <= 2'd0;
                txeq_done        <= 1'd0;
                end 
                
            //---------- Process TXEQ Preset ---------------
            2'd1    :
                begin
                fsm_tx           <= FSM_TXEQ_PRESET; 
                txeq_txcoeff     <= txeq_txcoeff;
                txeq_txcoeff_cnt <= 2'd0;
                txeq_done        <= 1'd0;
                end  
                
            //---------- Coefficient -----------------------
            2'd2    :
                begin
                fsm_tx           <= FSM_TXEQ_TXCOEFF; 
                txeq_txcoeff     <= {txeq_deemph_reg2, txeq_txcoeff[18:6]};
                txeq_txcoeff_cnt <= 2'd1;
                txeq_done        <= 1'd0;
                end
                
            //---------- Query -----------------------------
            2'd3    :
                begin
                fsm_tx           <= FSM_TXEQ_QUERY; 
                txeq_txcoeff     <= txeq_txcoeff;
                txeq_txcoeff_cnt <= 2'd0;
                txeq_done        <= 1'd0;
                end
                
            //---------- Default ---------------------------
            default :
                begin
                fsm_tx           <= FSM_TXEQ_IDLE; 
                txeq_txcoeff     <= txeq_txcoeff;
                txeq_txcoeff_cnt <= 2'd0;
                txeq_done        <= 1'd0;
                end
                
            endcase
            
            end
            
        //---------- Process TXEQ Preset -------------------
        FSM_TXEQ_PRESET :
        
            begin
            fsm_tx           <= (txeq_preset_done ? FSM_TXEQ_DONE : FSM_TXEQ_PRESET);
            txeq_txcoeff     <= txeq_preset;
            txeq_txcoeff_cnt <= 2'd0;
            txeq_done        <= 1'd0;
            end    
            
        //---------- Latch Link Partner TX Coefficient -----
        FSM_TXEQ_TXCOEFF :
        
            begin
            fsm_tx <= ((txeq_txcoeff_cnt == 2'd2) ? FSM_TXEQ_REMAP : FSM_TXEQ_TXCOEFF);
            
            //---------- Shift in extra bit for TXMAINCURSOR 
            if (txeq_txcoeff_cnt == 2'd1)
                txeq_txcoeff <= {1'd0, txeq_deemph_reg2, txeq_txcoeff[18:7]};
            else
                txeq_txcoeff <= {txeq_deemph_reg2, txeq_txcoeff[18:6]};
                
            txeq_txcoeff_cnt <= txeq_txcoeff_cnt + 2'd1;
            txeq_done        <= 1'd0; 
            end
            
        //---------- Remap to GT TX Coefficient ------------
        FSM_TXEQ_REMAP :
        
            begin
            fsm_tx           <= FSM_TXEQ_DONE;
            txeq_txcoeff     <= txeq_txcoeff << 1;          // Multiply by 2x
            txeq_txcoeff_cnt <= 2'd0;
            txeq_done        <= 1'd0; 
            end
            
        //---------- Query TXEQ Coefficient ----------------
        FSM_TXEQ_QUERY:
        
            begin
            fsm_tx           <= FSM_TXEQ_DONE;
            txeq_txcoeff     <= txeq_txcoeff; 
            txeq_txcoeff_cnt <= 2'd0;
            txeq_done        <= 1'd0;
            end     
                  
        //---------- Done ----------------------------------
        FSM_TXEQ_DONE :
        
            begin
            fsm_tx           <= ((txeq_control_reg2 == 2'd0) ? FSM_TXEQ_IDLE : FSM_TXEQ_DONE);
            txeq_txcoeff     <= txeq_txcoeff;          
            txeq_txcoeff_cnt <= 2'd0;
            txeq_done        <= 1'd1;
            end        
                          
        //---------- Default State -------------------------
        default : 
            begin
            fsm_tx           <=  FSM_TXEQ_IDLE;
            txeq_txcoeff     <= 19'd0;
            txeq_txcoeff_cnt <=  2'd0;
            txeq_done        <=  1'd0;
            end    
                    
        endcase
        
        end
        
end  



//---------- RXEQ FSM ----------------------------------------------------------
always @ (posedge EQ_CLK)
begin

    if (!EQ_RST_N)
        begin
        fsm_rx               <= FSM_RXEQ_IDLE; 
        rxeq_preset          <=  3'd0;
        rxeq_preset_valid    <=  1'd0;
        rxeq_txpreset        <=  4'd0;
        rxeq_txcoeff         <= 18'd0; 
        rxeq_cnt             <=  3'd0;
        rxeq_fs              <=  6'd0;
        rxeq_lf              <=  6'd0;
        rxeq_new_txcoeff_req <=  1'd0; 
        rxeq_new_txcoeff     <= 18'd0;
        rxeq_lffs_sel        <=  1'd0;
        rxeq_adapt_done_reg  <=  1'd0;
        rxeq_adapt_done      <=  1'd0;   
        rxeq_done            <=  1'd0; 
        end                    
    else
        begin
        
        case (fsm_rx)
        
        //---------- Idle State ----------------------------
        FSM_RXEQ_IDLE :
        
            begin
            
            case (rxeq_control_reg2)
                
            //---------- Process RXEQ Preset ---------------
            2'd1 :
                begin
                fsm_rx               <= FSM_RXEQ_PRESET; 
                rxeq_preset          <= rxeq_preset_reg2;
                rxeq_preset_valid    <= 1'd0;
                rxeq_txpreset        <= rxeq_txpreset;
                rxeq_txcoeff         <= rxeq_txcoeff;
                rxeq_cnt             <= 3'd0;
                rxeq_fs              <= rxeq_fs;
                rxeq_lf              <= rxeq_lf;
                rxeq_new_txcoeff_req <= 1'd0;
                rxeq_new_txcoeff     <= rxeq_new_txcoeff;
                rxeq_lffs_sel        <= 1'd0;
                rxeq_adapt_done_reg  <= 1'd0;
                rxeq_adapt_done      <= 1'd0;
                rxeq_done            <= 1'd0; 
                end  
                
            //---------- Request New TX Coefficient --------
            2'd2 :
                begin
                fsm_rx               <= FSM_RXEQ_TXCOEFF; 
                rxeq_preset          <= rxeq_preset;
                rxeq_preset_valid    <= 1'd0;
                rxeq_txpreset        <= rxeq_txpreset_reg2;
                rxeq_txcoeff         <= {txeq_deemph_reg2, rxeq_txcoeff[17:6]};
                rxeq_cnt             <= 3'd1;
                rxeq_fs              <= rxeq_lffs_reg2;
                rxeq_lf              <= rxeq_lf;
                rxeq_new_txcoeff_req <= 1'd0;
                rxeq_new_txcoeff     <= rxeq_new_txcoeff;
                rxeq_lffs_sel        <= 1'd0;
                rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
                rxeq_adapt_done      <= 1'd0;
                rxeq_done            <= 1'd0; 
                end
                
            //---------- Phase2/3 Bypass (reuse logic from rxeq_control = 2 ----
            2'd3 :
                begin
                fsm_rx               <= FSM_RXEQ_TXCOEFF; 
                rxeq_preset          <= rxeq_preset;
                rxeq_preset_valid    <= 1'd0;
                rxeq_txpreset        <= rxeq_txpreset_reg2;
                rxeq_txcoeff         <= {txeq_deemph_reg2, rxeq_txcoeff[17:6]};
                rxeq_cnt             <= 3'd1;
                rxeq_fs              <= rxeq_lffs_reg2;
                rxeq_lf              <= rxeq_lf;
                rxeq_new_txcoeff_req <= 1'd0;
                rxeq_new_txcoeff     <= rxeq_new_txcoeff;
                rxeq_lffs_sel        <= 1'd0;
                rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
                rxeq_adapt_done      <= 1'd0;
                rxeq_done            <= 1'd0; 
                end
                
            //---------- Default ---------------------------
            default :
                begin
                fsm_rx               <= FSM_RXEQ_IDLE; 
                rxeq_preset          <= rxeq_preset;
                rxeq_preset_valid    <= 1'd0;
                rxeq_txpreset        <= rxeq_txpreset;
                rxeq_txcoeff         <= rxeq_txcoeff;
                rxeq_cnt             <= 3'd0;
                rxeq_fs              <= rxeq_fs;
                rxeq_lf              <= rxeq_lf;
                rxeq_new_txcoeff_req <= 1'd0;
                rxeq_new_txcoeff     <= rxeq_new_txcoeff;
                rxeq_lffs_sel        <= 1'd0;
                rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
                rxeq_adapt_done      <= 1'd0;
                rxeq_done            <= 1'd0; 
                end
                
            endcase
            
            end
            
        //---------- Process RXEQ Preset -------------------
        FSM_RXEQ_PRESET :
        
            begin
            fsm_rx               <= (rxeqscan_preset_done ? FSM_RXEQ_DONE : FSM_RXEQ_PRESET);
            rxeq_preset          <= rxeq_preset_reg2;
            rxeq_preset_valid    <= 1'd1; 
            rxeq_txpreset        <= rxeq_txpreset;
            rxeq_txcoeff         <= rxeq_txcoeff; 
            rxeq_cnt             <= 3'd0;
            rxeq_fs              <= rxeq_fs;
            rxeq_lf              <= rxeq_lf;
            rxeq_new_txcoeff_req <= 1'd0;
            rxeq_new_txcoeff     <= rxeq_new_txcoeff;
            rxeq_lffs_sel        <= 1'd0;
            rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
            rxeq_adapt_done      <= 1'd0;
            rxeq_done            <= 1'd0; 
            end    
            
        //---------- Shift-in Link Partner TX Coefficient and Preset 
        FSM_RXEQ_TXCOEFF :
        
            begin
            fsm_rx               <= ((rxeq_cnt == 3'd2) ? FSM_RXEQ_LF : FSM_RXEQ_TXCOEFF);
            rxeq_preset          <= rxeq_preset;
            rxeq_preset_valid    <= 1'd0; 
            rxeq_txpreset        <= rxeq_txpreset_reg2;
            rxeq_txcoeff         <= {txeq_deemph_reg2, rxeq_txcoeff[17:6]}; 
            rxeq_cnt             <= rxeq_cnt + 2'd1;
            rxeq_fs              <= rxeq_fs;
            rxeq_lf              <= rxeq_lf;
            rxeq_new_txcoeff_req <= 1'd0;
            rxeq_new_txcoeff     <= rxeq_new_txcoeff;
            rxeq_lffs_sel        <= 1'd1;
            rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
            rxeq_adapt_done      <= 1'd0;
            rxeq_done            <= 1'd0; 
            end
            
        //---------- Read Low Frequency (LF) Value ---------
        FSM_RXEQ_LF :
            begin
            fsm_rx               <= ((rxeq_cnt == 3'd7) ? FSM_RXEQ_NEW_TXCOEFF_REQ : FSM_RXEQ_LF);
            rxeq_preset          <= rxeq_preset;
            rxeq_preset_valid    <= 1'd0; 
            rxeq_txpreset        <= rxeq_txpreset;
            rxeq_txcoeff         <= rxeq_txcoeff; 
            rxeq_cnt             <= rxeq_cnt + 2'd1;
            rxeq_fs              <= rxeq_fs;
            rxeq_lf              <= ((rxeq_cnt == 3'd7) ? rxeq_lffs_reg2 : rxeq_lf);
            rxeq_new_txcoeff_req <= 1'd0;
            rxeq_new_txcoeff     <= rxeq_new_txcoeff;
            rxeq_lffs_sel        <= 1'd1;
            rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
            rxeq_adapt_done      <= 1'd0;
            rxeq_done            <= 1'd0; 
            end
            
        //---------- Request New TX Coefficient ------------
        FSM_RXEQ_NEW_TXCOEFF_REQ :
        
            begin            
            rxeq_preset          <= rxeq_preset;
            rxeq_preset_valid    <= 1'd0; 
            rxeq_txpreset        <= rxeq_txpreset;
            rxeq_txcoeff         <= rxeq_txcoeff; 
            rxeq_cnt             <= 3'd0;
            rxeq_fs              <= rxeq_fs;
            rxeq_lf              <= rxeq_lf;
            
            if (rxeqscan_new_txcoeff_done)
                begin
                fsm_rx               <= FSM_RXEQ_DONE;
                rxeq_new_txcoeff_req <= 1'd0;
                rxeq_new_txcoeff     <= rxeqscan_lffs_sel ? {14'd0, rxeqscan_new_txcoeff[3:0]} : rxeqscan_new_txcoeff;
                rxeq_lffs_sel        <= rxeqscan_lffs_sel;
                rxeq_adapt_done_reg  <= rxeqscan_adapt_done || rxeq_adapt_done_reg;
                rxeq_adapt_done      <= rxeqscan_adapt_done || rxeq_adapt_done_reg;
                rxeq_done            <= 1'd1; 
                end
            else
                begin
                fsm_rx               <= FSM_RXEQ_NEW_TXCOEFF_REQ;
                rxeq_new_txcoeff_req <= 1'd1;
                rxeq_new_txcoeff     <= rxeq_new_txcoeff;
                rxeq_lffs_sel        <= 1'd0;
                rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
                rxeq_adapt_done      <= 1'd0;
                rxeq_done            <= 1'd0; 
                end
            
            end     
             
        //---------- RXEQ Done -----------------------------
        FSM_RXEQ_DONE :
        
            begin
            fsm_rx               <= ((rxeq_control_reg2 == 2'd0) ? FSM_RXEQ_IDLE : FSM_RXEQ_DONE);
            rxeq_preset          <= rxeq_preset;
            rxeq_preset_valid    <= 1'd0;
            rxeq_txpreset        <= rxeq_txpreset; 
            rxeq_txcoeff         <= rxeq_txcoeff;
            rxeq_cnt             <= 3'd0;
            rxeq_fs              <= rxeq_fs;
            rxeq_lf              <= rxeq_lf;
            rxeq_new_txcoeff_req <= 1'd0;
            rxeq_new_txcoeff     <= rxeq_new_txcoeff;
            rxeq_lffs_sel        <= rxeq_lffs_sel;
            rxeq_adapt_done_reg  <= rxeq_adapt_done_reg;
            rxeq_adapt_done      <= rxeq_adapt_done;  
            rxeq_done            <= 1'd1; 
            end        
                          
        //---------- Default State -------------------------
        default : 
            begin
            fsm_rx               <= FSM_RXEQ_IDLE;
            rxeq_preset          <=  3'd0;
            rxeq_preset_valid    <=  1'd0;
            rxeq_txpreset        <=  4'd0;
            rxeq_txcoeff         <= 18'd0;
            rxeq_cnt             <=  3'd0;
            rxeq_fs              <=  6'd0;
            rxeq_lf              <=  6'd0;
            rxeq_new_txcoeff_req <=  1'd0;
            rxeq_new_txcoeff     <= 18'd0;
            rxeq_lffs_sel        <=  1'd0;
            rxeq_adapt_done_reg  <=  1'd0;
            rxeq_adapt_done      <=  1'd0;
            rxeq_done            <=  1'd0;   
            end    
                    
    	   endcase
        
        end
        
end      



//---------- RXEQ Eye Scan Module ----------------------------------------------
model_ap2_tst_rxeq_scan #
(
    .PCIE_SIM_MODE                      (PCIE_SIM_MODE),
    .PCIE_GT_DEVICE                     (PCIE_GT_DEVICE),
    .PCIE_RXEQ_MODE_GEN3                (PCIE_RXEQ_MODE_GEN3)
)

model_ap2_tst_rxeq_scan_i
(

    //---------- Input -------------------------------------
    .RXEQSCAN_CLK                       (EQ_CLK),
    .RXEQSCAN_RST_N                     (EQ_RST_N),
    .RXEQSCAN_CONTROL                   (rxeq_control_reg2),
    .RXEQSCAN_FS                        (rxeq_fs),      
    .RXEQSCAN_LF                        (rxeq_lf), 
    .RXEQSCAN_PRESET                    (rxeq_preset),
    .RXEQSCAN_PRESET_VALID              (rxeq_preset_valid),   
    .RXEQSCAN_TXPRESET                  (rxeq_txpreset),
    .RXEQSCAN_TXCOEFF                   (rxeq_txcoeff),    
    .RXEQSCAN_NEW_TXCOEFF_REQ           (rxeq_new_txcoeff_req),                
    
    //---------- Output ------------------------------------
    .RXEQSCAN_PRESET_DONE               (rxeqscan_preset_done),
    .RXEQSCAN_NEW_TXCOEFF               (rxeqscan_new_txcoeff),
    .RXEQSCAN_NEW_TXCOEFF_DONE          (rxeqscan_new_txcoeff_done),
    .RXEQSCAN_LFFS_SEL                  (rxeqscan_lffs_sel),
    .RXEQSCAN_ADAPT_DONE                (rxeqscan_adapt_done)
    
); 



//---------- PIPE EQ Output ----------------------------------------------------
assign EQ_TXEQ_DEEMPH      = txeq_txcoeff[0];       
assign EQ_TXEQ_PRECURSOR   = gen3_reg2 ? txeq_txcoeff[ 4: 0] : 5'h00;
assign EQ_TXEQ_MAINCURSOR  = gen3_reg2 ? txeq_txcoeff[12: 6] : 7'h00; 
assign EQ_TXEQ_POSTCURSOR  = gen3_reg2 ? txeq_txcoeff[17:13] : 5'h00;
assign EQ_TXEQ_DEEMPH_OUT  = {1'd0, txeq_txcoeff[18:14], txeq_txcoeff[12:7], 1'd0, txeq_txcoeff[5:1]}; // Divide by 2x
assign EQ_TXEQ_DONE        = txeq_done;
assign EQ_TXEQ_FSM         = fsm_tx;

assign EQ_RXEQ_NEW_TXCOEFF = rxeq_user_en_reg2 ? rxeq_user_txcoeff_reg2 : rxeq_new_txcoeff;
assign EQ_RXEQ_LFFS_SEL    = rxeq_user_en_reg2 ? rxeq_user_mode_reg2    : rxeq_lffs_sel;
assign EQ_RXEQ_ADAPT_DONE  = rxeq_adapt_done;
assign EQ_RXEQ_DONE        = rxeq_done;
assign EQ_RXEQ_FSM         = fsm_rx;



endmodule



`timescale 1ns/1ps
module model_ap2_tst_rxeq_scan #
(

    parameter PCIE_SIM_MODE       = "FALSE",                // PCIe sim mode 
    parameter PCIE_GT_DEVICE      = "GTX",                  // PCIe GT device
    parameter PCIE_RXEQ_MODE_GEN3 = 1,                      // PCIe RX equalization mode
    parameter CONVERGE_MAX        = 22'd3125000,            // Convergence max count (12ms) 
    parameter CONVERGE_MAX_BYPASS = 22'd2083333             // Convergence max count for phase2/3 bypass mode (8ms)
)

(

    //---------- Input -------------------------------------
    input               RXEQSCAN_CLK,                      
    input               RXEQSCAN_RST_N,
       
    input       [ 1:0]  RXEQSCAN_CONTROL,   
    input       [ 2:0]  RXEQSCAN_PRESET,
    input               RXEQSCAN_PRESET_VALID,
    input       [ 3:0]  RXEQSCAN_TXPRESET,
    input       [17:0]  RXEQSCAN_TXCOEFF,
    input               RXEQSCAN_NEW_TXCOEFF_REQ,
    input       [ 5:0]  RXEQSCAN_FS,
    input       [ 5:0]  RXEQSCAN_LF,
     
    
    //---------- Output ------------------------------------
    output              RXEQSCAN_PRESET_DONE,
    output      [17:0]  RXEQSCAN_NEW_TXCOEFF,
    output              RXEQSCAN_NEW_TXCOEFF_DONE,
    output              RXEQSCAN_LFFS_SEL,
    output              RXEQSCAN_ADAPT_DONE

);

    //---------- Input Register ----------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 2:0]  preset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 preset_valid_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 3:0]  txpreset_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [17:0]  txcoeff_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 new_txcoeff_req_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  fs_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  lf_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 2:0]  preset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 preset_valid_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 3:0]  txpreset_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [17:0]  txcoeff_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 new_txcoeff_req_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  fs_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [ 5:0]  lf_reg2;

    //---------- Internal Signals --------------------------
    reg                 adapt_done_cnt = 1'd0;

    //---------- Output Register ---------------------------          
    reg                 preset_done      =  1'd0;
    reg         [21:0]  converge_cnt     = 22'd0;
    reg         [17:0]  new_txcoeff      = 18'd0;
    reg                 new_txcoeff_done =  1'd0;
    reg                 lffs_sel         =  1'd0;
    reg                 adapt_done       =  1'd0;
    reg         [ 3:0]  fsm              =  4'd0;

    //---------- FSM ---------------------------------------                                         
    localparam          FSM_IDLE            = 4'b0001;
    localparam          FSM_PRESET          = 4'b0010;
    localparam          FSM_CONVERGE        = 4'b0100;
    localparam          FSM_NEW_TXCOEFF_REQ = 4'b1000; 
    
    //---------- Simulation Speedup ------------------------
    //  Gen3:  32 bits / PCLK : 1 million bits / X PCLK
    //         X = 
    //------------------------------------------------------
    localparam converge_max_cnt        = (PCIE_SIM_MODE == "TRUE") ? 22'd1000 : CONVERGE_MAX;   
    localparam converge_max_bypass_cnt = (PCIE_SIM_MODE == "TRUE") ? 22'd1000 : CONVERGE_MAX_BYPASS;   
    
    

//---------- Input FF ----------------------------------------------------------
always @ (posedge RXEQSCAN_CLK)
begin

    if (!RXEQSCAN_RST_N)
        begin   
        //---------- 1st Stage FF --------------------------  
        preset_reg1          <=  3'd0;
        preset_valid_reg1    <=  1'd0;
        txpreset_reg1        <=  4'd0;
        txcoeff_reg1         <= 18'd0;
        new_txcoeff_req_reg1 <=  1'd0;
        fs_reg1              <=  6'd0;
        lf_reg1              <=  6'd0;
        //---------- 2nd Stage FF --------------------------
        preset_reg2          <=  3'd0;
        preset_valid_reg2    <=  1'd0;
        txpreset_reg2        <=  4'd0;
        txcoeff_reg2         <= 18'd0;
        new_txcoeff_req_reg2 <=  1'd0;
        fs_reg2              <=  6'd0;
        lf_reg2              <=  6'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------  
        preset_reg1          <= RXEQSCAN_PRESET;
        preset_valid_reg1    <= RXEQSCAN_PRESET_VALID;
        txpreset_reg1        <= RXEQSCAN_TXPRESET;
        txcoeff_reg1         <= RXEQSCAN_TXCOEFF;
        new_txcoeff_req_reg1 <= RXEQSCAN_NEW_TXCOEFF_REQ;
        fs_reg1              <= RXEQSCAN_FS;
        lf_reg1              <= RXEQSCAN_LF;
        //---------- 2nd Stage FF -------------------------- 
        preset_reg2          <= preset_reg1;
        preset_valid_reg2    <= preset_valid_reg1;
        txpreset_reg2        <= txpreset_reg1;
        txcoeff_reg2         <= txcoeff_reg1;
        new_txcoeff_req_reg2 <= new_txcoeff_req_reg1;
        fs_reg2              <= fs_reg1;
        lf_reg2              <= lf_reg1;
        end
        
end     



//---------- Eye Scan ----------------------------------------------------------
always @ (posedge RXEQSCAN_CLK)
begin

    if (!RXEQSCAN_RST_N)
        begin
        fsm              <=  FSM_IDLE;
        preset_done      <=  1'd0;
        converge_cnt     <= 22'd0;
        new_txcoeff      <= 18'd0;
        new_txcoeff_done <=  1'd0;
        lffs_sel         <=  1'd0;
        adapt_done       <=  1'd0;
        adapt_done_cnt   <=  1'd0;
        end                   
    else
    
        begin
    
        case (fsm)
        
        //---------- Idle State ----------------------------
        FSM_IDLE : 
            
            begin   
             
            //---------- Process RXEQ Preset ---------------
            if (preset_valid_reg2)
                begin
                fsm              <=  FSM_PRESET;
                preset_done      <=  1'd1;
                converge_cnt     <= 22'd0;
                new_txcoeff      <=  new_txcoeff;
                new_txcoeff_done <=  1'd0;
                lffs_sel         <=  1'd0;
                adapt_done       <=  1'd0;
                adapt_done_cnt   <=  adapt_done_cnt;
                end            
            //---------- Request New TX Coefficient --------
            else if (new_txcoeff_req_reg2)
                begin
                fsm              <=  FSM_CONVERGE;
                preset_done      <=  1'd0;
                converge_cnt     <= 22'd0;
              //new_txcoeff      <= (PCIE_RXEQ_MODE_GEN3 == 0) ? txcoeff_reg2 : 18'd4;  // Default
                new_txcoeff      <= (PCIE_RXEQ_MODE_GEN3 == 0) ? txcoeff_reg2 : (PCIE_GT_DEVICE == "GTX") ? 18'd5 : 18'd4;  // Optimized for Gen3 RX JTOL
                new_txcoeff_done <=  1'd0;
                lffs_sel         <= (PCIE_RXEQ_MODE_GEN3 == 0) ? 1'd0 : 1'd1;
                adapt_done       <=  1'd0; 
                adapt_done_cnt   <=  adapt_done_cnt;
                end  
            //---------- Default ---------------------------
            else
                begin
                fsm              <=  FSM_IDLE;
                preset_done      <=  1'd0;
                converge_cnt     <= 22'd0;
                new_txcoeff      <=  new_txcoeff;
                new_txcoeff_done <=  1'd0;
                lffs_sel         <=  1'd0;
                adapt_done       <=  1'd0;
                adapt_done_cnt   <=  adapt_done_cnt;
                end
                
            end
            
        //---------- Process RXEQ Preset -------------------
        FSM_PRESET :

            begin
            fsm              <= (!preset_valid_reg2) ? FSM_IDLE : FSM_PRESET;
            preset_done      <=  1'd1;
            converge_cnt     <= 22'd0;
            new_txcoeff      <=  new_txcoeff;
            new_txcoeff_done <=  1'd0;
            lffs_sel         <=  1'd0;
            adapt_done       <=  1'd0;
            adapt_done_cnt   <=  adapt_done_cnt;
            end
            
        //---------- Wait for Convergence ------------------    
        FSM_CONVERGE :
           
            begin
            if ((adapt_done_cnt == 1'd0) && (RXEQSCAN_CONTROL == 2'd2))
                begin
                fsm              <= FSM_NEW_TXCOEFF_REQ;
                preset_done      <=  1'd0;
                converge_cnt     <= 22'd0;
                new_txcoeff      <= new_txcoeff;
                new_txcoeff_done <= 1'd0;
                lffs_sel         <= lffs_sel;
                adapt_done       <= 1'd0;
                adapt_done_cnt   <= adapt_done_cnt;
                end
            else
                begin
                
                //---------- Phase2/3 ----------------------
                if (RXEQSCAN_CONTROL == 2'd2)
                    fsm <= (converge_cnt == converge_max_cnt)        ? FSM_NEW_TXCOEFF_REQ : FSM_CONVERGE;
                //---------- Phase2/3 Bypass ---------------
                else
                    fsm <= (converge_cnt == converge_max_bypass_cnt) ? FSM_NEW_TXCOEFF_REQ : FSM_CONVERGE;
                
                preset_done      <= 1'd0;
                converge_cnt     <= converge_cnt + 1'd1;
                new_txcoeff      <= new_txcoeff;
                new_txcoeff_done <= 1'd0;
                lffs_sel         <= lffs_sel;
                adapt_done       <= 1'd0;
                adapt_done_cnt   <= adapt_done_cnt;
                end
            end
            
        //---------- Request New TX Coefficient ------------
        FSM_NEW_TXCOEFF_REQ :

            begin 
            if (!new_txcoeff_req_reg2)
                begin
                fsm              <= FSM_IDLE;
                preset_done      <=  1'd0;
                converge_cnt     <= 22'd0;
                new_txcoeff      <= new_txcoeff;
                new_txcoeff_done <= 1'd0;
                lffs_sel         <= lffs_sel;
                adapt_done       <= 1'd0;
                adapt_done_cnt   <= (RXEQSCAN_CONTROL == 2'd3) ? 1'd0 : adapt_done_cnt + 1'd1;
                end
            else
                begin
                fsm              <= FSM_NEW_TXCOEFF_REQ;
                preset_done      <=  1'd0;
                converge_cnt     <= 22'd0;
                new_txcoeff      <= new_txcoeff;
                new_txcoeff_done <= 1'd1;
                lffs_sel         <= lffs_sel;
                adapt_done       <= (adapt_done_cnt == 1'd1) || (RXEQSCAN_CONTROL == 2'd3);
                adapt_done_cnt   <= adapt_done_cnt;
                end
            end
            
        //---------- Default State -------------------------
        default :
        
            begin
            fsm              <=  FSM_IDLE;
            preset_done      <=  1'd0;
            converge_cnt     <= 22'd0;
            new_txcoeff      <= 18'd0;
            new_txcoeff_done <=  1'd0;
            lffs_sel         <=  1'd0;
            adapt_done       <=  1'd0;
            adapt_done_cnt   <=  1'd0;
            end    

        endcase
        
        end
        
end



//---------- RXEQ Eye Scan Output ----------------------------------------------
assign RXEQSCAN_PRESET_DONE      = preset_done;     
assign RXEQSCAN_NEW_TXCOEFF      = new_txcoeff;
assign RXEQSCAN_NEW_TXCOEFF_DONE = new_txcoeff_done; 
assign RXEQSCAN_LFFS_SEL         = lffs_sel;  
assign RXEQSCAN_ADAPT_DONE       = adapt_done;



endmodule



`timescale 1ns/1ps
module model_ap2_tst_gt_common #(

parameter PCIE_SIM_MODE    = "FALSE",   // PCIe sim mode
parameter PCIE_GT_DEVICE   = "GTX",     // PCIe GT device
parameter PCIE_USE_MODE    = "2.1",     // PCIe use mode
parameter PCIE_PLL_SEL     = "CPLL",    // PCIe PLL select for Gen1/Gen2 only
parameter PCIE_REFCLK_FREQ = 0          // PCIe reference clock frequency
)

(
input                   CPLLPDREFCLK,
input               	PIPE_CLK,
input               	QPLL_QPLLPD,
input               	QPLL_QPLLRESET,
input               	QPLL_DRP_CLK,
input               	QPLL_DRP_RST_N,
input               	QPLL_DRP_OVRD,
input               	QPLL_DRP_GEN3,
input               	QPLL_DRP_START,
output      [5:0]  	QPLL_DRP_CRSCODE,
output      [8:0]  	QPLL_DRP_FSM,
output                  QPLL_DRP_DONE,
output                  QPLL_DRP_RESET,
output                  QPLL_QPLLLOCK,
output                  QPLL_QPLLOUTCLK,
output                  QPLL_QPLLOUTREFCLK
);

    //---------- QPLL DRP Module Output --------------------

wire        [7:0]  qpll_drp_addr;
wire               qpll_drp_en;
wire        [15:0] qpll_drp_di;
wire               qpll_drp_we;

   //---------- QPLL Wrapper Output -----------------------

wire        [15:0] qpll_drp_do;
wire               qpll_drp_rdy;

   //---------- QPLL Resets -----------------------


        //---------- QPLL DRP Module ---------------------------------------

model_ap2_tst_qpll_drp #
        (

	        .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),               // PCIe GT device
	        .PCIE_USE_MODE                  (PCIE_USE_MODE),                // PCIe use mode
	        .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                 // PCIe PLL select for Gen1/Gen2 only
	        .PCIE_REFCLK_FREQ               (PCIE_REFCLK_FREQ)              // PCIe reference clock frequency

        )
        model_ap2_tst_qpll_drp_i
        (

        //---------- Input -------------------------
	    .DRP_CLK                        (QPLL_DRP_CLK),
            .DRP_RST_N                      (!QPLL_DRP_RST_N),
            .DRP_OVRD                       (QPLL_DRP_OVRD),
            .DRP_GEN3                       (&QPLL_DRP_GEN3),
            .DRP_QPLLLOCK                   (QPLL_QPLLLOCK),
            .DRP_START                      (QPLL_DRP_START),
            .DRP_DO                         (qpll_drp_do),
            .DRP_RDY                        (qpll_drp_rdy),
																													     
        //----------           Output ------------------------
            .DRP_ADDR                       (qpll_drp_addr),
            .DRP_EN                         (qpll_drp_en),
            .DRP_DI                         (qpll_drp_di),
            .DRP_WE                         (qpll_drp_we),
            .DRP_DONE                       (QPLL_DRP_DONE),
            .DRP_QPLLRESET                  (QPLL_DRP_RESET),
            .DRP_CRSCODE                    (QPLL_DRP_CRSCODE),
            .DRP_FSM                        (QPLL_DRP_FSM)
        );


        //---------- QPLL Wrapper ------------------------------------------
model_ap2_tst_qpll_wrapper #
        (
	        .PCIE_SIM_MODE                  (PCIE_SIM_MODE),                // PCIe sim mode
	        .PCIE_GT_DEVICE                 (PCIE_GT_DEVICE),               // PCIe GT device
	        .PCIE_USE_MODE                  (PCIE_USE_MODE),                // PCIe use mode
	        .PCIE_PLL_SEL                   (PCIE_PLL_SEL),                 // PCIe PLL select for Gen1/Gen2 only
	        .PCIE_REFCLK_FREQ               (PCIE_REFCLK_FREQ)              // PCIe reference clock frequency
        )
        model_ap2_tst_qpll_wrapper_i
        (
        //---------- QPLL Clock Ports --------------
            .QPLL_CPLLPDREFCLK              (CPLLPDREFCLK),
            .QPLL_GTGREFCLK                 (PIPE_CLK),
            .QPLL_QPLLLOCKDETCLK            (1'd0),
            .QPLL_QPLLOUTCLK                (QPLL_QPLLOUTCLK),
            .QPLL_QPLLOUTREFCLK             (QPLL_QPLLOUTREFCLK),
            .QPLL_QPLLLOCK                  (QPLL_QPLLLOCK),
        //---------- QPLL Reset Ports --------------
            .QPLL_QPLLPD                    (QPLL_QPLLPD),
            .QPLL_QPLLRESET                 (QPLL_QPLLRESET),
        //---------- QPLL DRP Ports ----------------
            .QPLL_DRPCLK                    (QPLL_DRP_CLK),
            .QPLL_DRPADDR                   (qpll_drp_addr),
            .QPLL_DRPEN                     (qpll_drp_en),
            .QPLL_DRPDI                     (qpll_drp_di),
            .QPLL_DRPWE                     (qpll_drp_we),
            .QPLL_DRPDO                     (qpll_drp_do),
            .QPLL_DRPRDY                    (qpll_drp_rdy)			
        );
  
endmodule



`timescale 1ns/1ps
module model_ap2_tst_qpll_drp #
(

    parameter PCIE_GT_DEVICE   = "GTX",                     // PCIe GT device
    parameter PCIE_USE_MODE    = "3.0",                     // PCIe use mode
    parameter PCIE_PLL_SEL     = "CPLL",                    // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_REFCLK_FREQ = 0,                         // PCIe reference clock frequency
    parameter LOAD_CNT_MAX     = 2'd3,                      // Load max count
    parameter INDEX_MAX        = 3'd6                       // Index max count
        
)

(
    
    //---------- Input -------------------------------------
    input               DRP_CLK,
    input               DRP_RST_N,
    input               DRP_OVRD,
    input               DRP_GEN3,
    input               DRP_QPLLLOCK,
    input               DRP_START,
    input       [15:0]  DRP_DO,
    input               DRP_RDY,
    
    //---------- Output ------------------------------------
    output      [ 7:0]  DRP_ADDR,
    output              DRP_EN,  
    output      [15:0]  DRP_DI,   
    output              DRP_WE,
    output              DRP_DONE,
    output              DRP_QPLLRESET,
    output      [ 5:0]  DRP_CRSCODE,
    output      [ 8:0]  DRP_FSM
    
);

    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 ovrd_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 qplllock_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg1;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg1;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 ovrd_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 gen3_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 qplllock_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 start_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [15:0]  do_reg2;
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                 rdy_reg2;
    
    //---------- Internal Signals --------------------------
    reg         [ 1:0]  load_cnt =  2'd0;
    reg         [ 2:0]  index    =  3'd0;
    reg                 mode     =  1'd0;
    reg         [ 5:0]  crscode  =  6'd0;
    
    //---------- Output Registers --------------------------
    reg         [ 7:0]  addr    =  8'd0;
    reg         [15:0]  di      = 16'd0;
    reg                 done    =  1'd0;
    reg         [ 8:0]  fsm     =  7'd1;      
                        
    //---------- DRP Address -------------------------------  
    localparam          ADDR_QPLL_FBDIV               = 8'h36;
    localparam          ADDR_QPLL_CFG                 = 8'h32;
    localparam          ADDR_QPLL_LPF                 = 8'h31;  
    localparam          ADDR_CRSCODE                  = 8'h88;  
    localparam          ADDR_QPLL_COARSE_FREQ_OVRD    = 8'h35;
    localparam          ADDR_QPLL_COARSE_FREQ_OVRD_EN = 8'h36;  
    localparam          ADDR_QPLL_LOCK_CFG            = 8'h34;
    
    //---------- DRP Mask ----------------------------------
    localparam          MASK_QPLL_FBDIV               = 16'b1111110000000000;  // Unmask bit [ 9: 0] 
    localparam          MASK_QPLL_CFG                 = 16'b1111111110111111;  // Unmask bit [    6]
    localparam          MASK_QPLL_LPF                 = 16'b1000011111111111;  // Unmask bit [14:11]
    localparam          MASK_QPLL_COARSE_FREQ_OVRD    = 16'b0000001111111111;  // Unmask bit [15:10] 
    localparam          MASK_QPLL_COARSE_FREQ_OVRD_EN = 16'b1111011111111111;  // Unmask bit [   11]      
    localparam          MASK_QPLL_LOCK_CFG            = 16'b1110011111111111;  // Unmask bit [12:11]     

    //---------- DRP Data for Normal QPLLLOCK Mode ---------
    localparam          NORM_QPLL_COARSE_FREQ_OVRD    = 16'b0000000000000000;  // Coarse freq value
    localparam          NORM_QPLL_COARSE_FREQ_OVRD_EN = 16'b0000000000000000;  // Normal QPLL lock  
    localparam          NORM_QPLL_LOCK_CFG            = 16'b0000000000000000;  // Normal QPLL lock config 
     
    //---------- DRP Data for Optimize QPLLLOCK Mode -------
    localparam          OVRD_QPLL_COARSE_FREQ_OVRD    = 16'b0000000000000000;  // Coarse freq value
    localparam          OVRD_QPLL_COARSE_FREQ_OVRD_EN = 16'b0000100000000000;  // Override QPLL lock 
    localparam          OVRD_QPLL_LOCK_CFG            = 16'b0000000000000000;  // Override QPLL lock config 
    
    //---------- Select QPLL Feedback Divider --------------
    //  N = 100 for 100 MHz ref clk and 10Gb/s line rate
    //  N =  80 for 125 MHz ref clk and 10Gb/s line rate
    //  N =  40 for 250 MHz ref clk and 10Gb/s line rate
    //------------------------------------------------------
    //  N =  80 for 100 MHz ref clk and  8Gb/s line rate
    //  N =  64 for 125 MHz ref clk and  8Gb/s line rate
    //  N =  32 for 250 MHz ref clk and  8Gb/s line rate
    //------------------------------------------------------
    localparam          QPLL_FBDIV = (PCIE_REFCLK_FREQ == 2) && (PCIE_PLL_SEL == "QPLL") ? 16'b0000000010000000 : 
                                     (PCIE_REFCLK_FREQ == 1) && (PCIE_PLL_SEL == "QPLL") ? 16'b0000000100100000 : 
                                     (PCIE_REFCLK_FREQ == 0) && (PCIE_PLL_SEL == "QPLL") ? 16'b0000000101110000 : 
                                     (PCIE_REFCLK_FREQ == 2) && (PCIE_PLL_SEL == "CPLL") ? 16'b0000000001100000 : 
                                     (PCIE_REFCLK_FREQ == 1) && (PCIE_PLL_SEL == "CPLL") ? 16'b0000000011100000 : 16'b0000000100100000;
    
    localparam          GEN12_QPLL_FBDIV = (PCIE_REFCLK_FREQ == 2) ? 16'b0000000010000000 : 
                                           (PCIE_REFCLK_FREQ == 1) ? 16'b0000000100100000 : 16'b0000000101110000;

    localparam          GEN3_QPLL_FBDIV  = (PCIE_REFCLK_FREQ == 2) ? 16'b0000000001100000 : 
                                           (PCIE_REFCLK_FREQ == 1) ? 16'b0000000011100000 : 16'b0000000100100000;
     
    //---------- Select QPLL Configuration ---------------------------
    //  QPLL_CFG[6] = 0 for upper band
    //              = 1 for lower band
    //----------------------------------------------------------------
    localparam          GEN12_QPLL_CFG = (PCIE_PLL_SEL == "QPLL") ? 16'b0000000000000000 : 16'b0000000001000000;
    localparam          GEN3_QPLL_CFG  = 16'b0000000001000000;  
     
    //---------- Select QPLL LPF -------------------------------------
    localparam          GEN12_QPLL_LPF = (PCIE_PLL_SEL == "QPLL") ? 16'b0_0100_00000000000 : 16'b0_1101_00000000000;
    localparam          GEN3_QPLL_LPF  = 16'b0_1101_00000000000;  
     
     
     
    //---------- DRP Data ----------------------------------       
    wire        [15:0]  data_qpll_fbdiv;  
    wire        [15:0]  data_qpll_cfg;  
    wire        [15:0]  data_qpll_lpf;  
    wire        [15:0]  data_qpll_coarse_freq_ovrd;               
    wire        [15:0]  data_qpll_coarse_freq_ovrd_en; 
    wire        [15:0]  data_qpll_lock_cfg;      
           
    //---------- FSM ---------------------------------------  
    localparam          FSM_IDLE      = 9'b000000001;  
    localparam          FSM_LOAD      = 9'b000000010;                           
    localparam          FSM_READ      = 9'b000000100;
    localparam          FSM_RRDY      = 9'b000001000;
    localparam          FSM_WRITE     = 9'b000010000;
    localparam          FSM_WRDY      = 9'b000100000;    
    localparam          FSM_DONE      = 9'b001000000; 
    localparam          FSM_QPLLRESET = 9'b010000000; 
    localparam          FSM_QPLLLOCK  = 9'b100000000;


    
//---------- Input FF ----------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        //---------- 1st Stage FF --------------------------
        ovrd_reg1     <=  1'd0;
        gen3_reg1     <=  1'd0;
        qplllock_reg1 <=  1'd0;
        start_reg1    <=  1'd0;
        do_reg1       <= 16'd0;
        rdy_reg1      <=  1'd0;
        //---------- 2nd Stage FF --------------------------
        ovrd_reg2     <=  1'd0;
        gen3_reg2     <=  1'd0;
        qplllock_reg2 <=  1'd0;
        start_reg2    <=  1'd0;
        do_reg2       <= 16'd0;
        rdy_reg2      <=  1'd0;
        end
        
    else
        begin
        //---------- 1st Stage FF --------------------------
        ovrd_reg1     <= DRP_OVRD;
        gen3_reg1     <= DRP_GEN3;
        qplllock_reg1 <= DRP_QPLLLOCK;
        start_reg1    <= DRP_START;
        do_reg1       <= DRP_DO;
        rdy_reg1      <= DRP_RDY;
        //---------- 2nd Stage FF --------------------------
        ovrd_reg2     <= ovrd_reg1;
        gen3_reg2     <= gen3_reg1;
        qplllock_reg2 <= qplllock_reg1;
        start_reg2    <= start_reg1;
        do_reg2       <= do_reg1;
        rdy_reg2      <= rdy_reg1;
        end
    
end  



//---------- Select DRP Data ---------------------------------------------------
assign data_qpll_fbdiv               = (gen3_reg2) ? GEN3_QPLL_FBDIV : GEN12_QPLL_FBDIV;
assign data_qpll_cfg                 = (gen3_reg2) ? GEN3_QPLL_CFG   : GEN12_QPLL_CFG;
assign data_qpll_lpf                 = (gen3_reg2) ? GEN3_QPLL_LPF   : GEN12_QPLL_LPF;
assign data_qpll_coarse_freq_ovrd    =  NORM_QPLL_COARSE_FREQ_OVRD;
assign data_qpll_coarse_freq_ovrd_en = (ovrd_reg2) ? OVRD_QPLL_COARSE_FREQ_OVRD_EN : NORM_QPLL_COARSE_FREQ_OVRD_EN;
assign data_qpll_lock_cfg            = (ovrd_reg2) ? OVRD_QPLL_LOCK_CFG            : NORM_QPLL_LOCK_CFG;


//---------- Load Counter ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        load_cnt <= 2'd0;
    else
    
        //---------- Increment Load Counter ----------------
        if ((fsm == FSM_LOAD) && (load_cnt < LOAD_CNT_MAX))
            load_cnt <= load_cnt + 2'd1;
            
        //---------- Hold Load Counter ---------------------
        else if ((fsm == FSM_LOAD) && (load_cnt == LOAD_CNT_MAX))
            load_cnt <= load_cnt;
            
        //---------- Reset Load Counter --------------------
        else
            load_cnt <= 2'd0;
        
end 



//---------- Update DRP Address and Data ---------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        addr    <=  8'd0;
        di      <= 16'd0;
        crscode <=  6'd0;
        end
    else
        begin
        
        case (index)

        //--------------------------------------------------    
        3'd0 :
            begin        
            addr    <= ADDR_QPLL_FBDIV;
            di      <= (do_reg2 & MASK_QPLL_FBDIV) | (mode ? data_qpll_fbdiv : QPLL_FBDIV);
            crscode <= crscode;
            end   
                
        //--------------------------------------------------    
        3'd1 :
            begin       
            addr    <= ADDR_QPLL_CFG;
            if (PCIE_GT_DEVICE == "GTX") 
                di <= (do_reg2 & MASK_QPLL_CFG) | data_qpll_cfg;
            else
                di <= (do_reg2 & 16'hFFFF) | data_qpll_cfg;
            crscode <= crscode;
            end       
            
        //--------------------------------------------------    
        3'd2 :
            begin        
            addr    <= ADDR_QPLL_LPF;
            if (PCIE_GT_DEVICE == "GTX") 
                di <= (do_reg2 & MASK_QPLL_LPF) | data_qpll_lpf;
            else
                di <= (do_reg2 & 16'hFFFF) | data_qpll_lpf;
            crscode <= crscode;
            end     
                
        //--------------------------------------------------
        3'd3 :
            begin        
            addr <= ADDR_CRSCODE;
            di   <= do_reg2;
            
            //---------- Latch CRS Code --------------------
            if (ovrd_reg2)
                crscode <= do_reg2[6:1];                 
            else
                crscode <= crscode;   
            end
           
        //--------------------------------------------------    
        3'd4 :
            begin        
            addr    <= ADDR_QPLL_COARSE_FREQ_OVRD;
            di      <= (do_reg2 & MASK_QPLL_COARSE_FREQ_OVRD) | {(crscode - 6'd1), data_qpll_coarse_freq_ovrd[9:0]};
            crscode <= crscode;
            end    
            
        //--------------------------------------------------    
        3'd5 :
            begin        
            addr    <= ADDR_QPLL_COARSE_FREQ_OVRD_EN;
            di      <= (do_reg2 & MASK_QPLL_COARSE_FREQ_OVRD_EN) | data_qpll_coarse_freq_ovrd_en;
            crscode <= crscode;
            end    
            
        //--------------------------------------------------    
        3'd6 :
            begin        
            addr    <= ADDR_QPLL_LOCK_CFG;
            di      <= (do_reg2 & MASK_QPLL_LOCK_CFG) | data_qpll_lock_cfg;
            crscode <= crscode;
            end       
            
        //--------------------------------------------------
        default : 
            begin
            addr    <=  8'd0;
            di      <= 16'd0;
            crscode <=  6'd0;
            end
            
        endcase
        
        end
        
end  



//---------- QPLL DRP FSM ------------------------------------------------------
always @ (posedge DRP_CLK)
begin

    if (!DRP_RST_N)
        begin
        fsm   <= FSM_IDLE;
        index <= 3'd0;
        mode  <= 1'd0;
        done  <= 1'd0;
        end
    else
        begin
        
        case (fsm)

        //---------- Idle State ----------------------------
        FSM_IDLE :  
          
            begin
            if (start_reg2)
                begin
                fsm   <= FSM_LOAD;
                index <= 3'd0;
                mode  <= 1'd0;
                done  <= 1'd0;
                end
            else if ((gen3_reg2 != gen3_reg1) && (PCIE_PLL_SEL == "QPLL"))
                begin
                fsm   <= FSM_LOAD;
                index <= 3'd0;
                mode  <= 1'd1;
                done  <= 1'd0;
                end
            else
                begin
                fsm   <= FSM_IDLE;
                index <= 3'd0;
                mode  <= 1'd0;
                done  <= 1'd1;
                end
            end    
            
        //---------- Load DRP Address  ---------------------
        FSM_LOAD :
        
            begin
            fsm   <= (load_cnt == LOAD_CNT_MAX) ? FSM_READ : FSM_LOAD;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end  
            
        //---------- Read DRP ------------------------------
        FSM_READ :
        
            begin
            fsm   <= FSM_RRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end
            
        //---------- Read DRP Ready ------------------------
        FSM_RRDY :    
        
            begin
            fsm   <= (rdy_reg2 ? FSM_WRITE : FSM_RRDY);
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end  
            
        //---------- Write DRP -----------------------------
        FSM_WRITE :    
        
            begin
            fsm   <= FSM_WRDY;
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end       
            
        //---------- Write DRP Ready -----------------------
        FSM_WRDY :    
        
            begin
            fsm   <= (rdy_reg2 ? FSM_DONE : FSM_WRDY);
            index <= index;
            mode  <= mode;
            done  <= 1'd0;
            end        
             
        //---------- DRP Done ------------------------------
        FSM_DONE :
        
            begin
            if ((index == INDEX_MAX) || (mode && (index == 3'd2)))
                begin
                fsm   <= mode ? FSM_QPLLRESET : FSM_IDLE;
                index <= 3'd0;
                mode  <= mode;
                done  <= 1'd0;
                end
            else       
                begin
                fsm   <= FSM_LOAD;
                index <= index + 3'd1;
                mode  <= mode;
                done  <= 1'd0;
                end
            end     
        
        //---------- QPLL Reset ----------------------------      
        FSM_QPLLRESET :
        
            begin
            fsm   <= !qplllock_reg2 ? FSM_QPLLLOCK : FSM_QPLLRESET;
            index <= 3'd0;
            mode  <= mode;
            done  <= 1'd0;
            end
            
        //---------- QPLL Reset ----------------------------      
        FSM_QPLLLOCK :
        
            begin
            fsm   <= qplllock_reg2 ? FSM_IDLE : FSM_QPLLLOCK;
            index <= 3'd0;
            mode  <= mode;
            done  <= 1'd0;
            end
              
        //---------- Default State -------------------------
        default :
        
            begin      
            fsm   <= FSM_IDLE;
            index <= 3'd0;
            mode  <= 1'd0;
            done  <= 1'd0;
            end
            
        endcase
        
        end
        
end 



//---------- QPLL DRP Output ---------------------------------------------------
assign DRP_ADDR      = addr;
assign DRP_EN        = (fsm == FSM_READ) || (fsm == FSM_WRITE);
assign DRP_DI        = di;
assign DRP_WE        = (fsm == FSM_WRITE); // || (fsm == FSM_WRDY);
assign DRP_DONE      = done;
assign DRP_QPLLRESET = (fsm == FSM_QPLLRESET);
assign DRP_CRSCODE   = crscode;
assign DRP_FSM       = fsm;



endmodule



`timescale 1ns/1ps
module model_ap2_tst_qpll_wrapper #
(
    
    parameter PCIE_SIM_MODE    = "FALSE",                   // PCIe sim mode
    parameter PCIE_GT_DEVICE   = "GTX",                     // PCIe GT device
    parameter PCIE_USE_MODE    = "3.0",                     // PCIe use mode
    parameter PCIE_PLL_SEL     = "CPLL",                    // PCIe PLL select for Gen1/Gen2 only
    parameter PCIE_REFCLK_FREQ = 0                          // PCIe reference clock frequency
 
)

(    
    
    //---------- QPLL Clock Ports --------------------------
    input               QPLL_CPLLPDREFCLK,
    input               QPLL_GTGREFCLK,
    input               QPLL_QPLLLOCKDETCLK,
    
    output              QPLL_QPLLOUTCLK,
    output              QPLL_QPLLOUTREFCLK,
    output              QPLL_QPLLLOCK,
    
    //---------- QPLL Reset Ports --------------------------
    input               QPLL_QPLLPD,
    input               QPLL_QPLLRESET,

    //---------- QPLL DRP Ports ----------------------------
    input               QPLL_DRPCLK,
    input       [ 7:0]  QPLL_DRPADDR,
    input               QPLL_DRPEN,
    input       [15:0]  QPLL_DRPDI,
    input               QPLL_DRPWE,
    
    output      [15:0]  QPLL_DRPDO,
    output              QPLL_DRPRDY
    
);



    //---------- Select QPLL Feedback Divider --------------
    //  N = 100 for 100 MHz ref clk and 10Gb/s line rate
    //  N =  80 for 125 MHz ref clk and 10Gb/s line rate
    //  N =  40 for 250 MHz ref clk and 10Gb/s line rate
    //------------------------------------------------------
    //  N =  80 for 100 MHz ref clk and  8Gb/s line rate
    //  N =  64 for 125 MHz ref clk and  8Gb/s line rate
    //  N =  32 for 250 MHz ref clk and  8Gb/s line rate
    //------------------------------------------------------
    localparam QPLL_FBDIV = (PCIE_REFCLK_FREQ == 2) && (PCIE_PLL_SEL == "QPLL") ? 10'b0010000000 : 
                            (PCIE_REFCLK_FREQ == 1) && (PCIE_PLL_SEL == "QPLL") ? 10'b0100100000 : 
                            (PCIE_REFCLK_FREQ == 0) && (PCIE_PLL_SEL == "QPLL") ? 10'b0101110000 : 
                            (PCIE_REFCLK_FREQ == 2) && (PCIE_PLL_SEL == "CPLL") ? 10'b0001100000 : 
                            (PCIE_REFCLK_FREQ == 1) && (PCIE_PLL_SEL == "CPLL") ? 10'b0011100000 : 10'b0100100000;
    
    //---------- Select GTP QPLL Feedback Divider ----------                     
    localparam GTP_QPLL_FBDIV  = (PCIE_REFCLK_FREQ == 2) ? 3'd2 :
                                 (PCIE_REFCLK_FREQ == 1) ? 3'd4 : 3'd5;

    //---------- Select BIAS_CFG ---------------------------
    localparam BIAS_CFG = ((PCIE_USE_MODE == "1.0") && (PCIE_PLL_SEL == "CPLL")) ? 64'h0000042000001000 : 64'h0000040000001000;


    wire cpllpd;        
    wire cpllrst;       

//---------- Select GTX or GTH or GTP ------------------------------------------
//  Notes  :  Attributes that are commented out uses the GT default settings
//------------------------------------------------------------------------------
generate if (PCIE_GT_DEVICE == "GTP") 

    //---------- GTP Common ----------------------------------------------------
    begin : gtp_common

    //---------- GTP Common Module ---------------------------------------------
    GTPE2_COMMON #
    (
       
        //---------- Simulation Attributes -------------------------------------                                                     
        .SIM_PLL0REFCLK_SEL             (3'b001),                               //                                                   
        .SIM_PLL1REFCLK_SEL             (3'b001),                               //                                                   
        .SIM_RESET_SPEEDUP              (PCIE_SIM_MODE),                        //                                                   
        .SIM_VERSION                    (PCIE_USE_MODE),                        //                                                   
                                                                                                                                     
        //---------- Clock Attributes ------------------------------------------                                                     
        .PLL0_CFG                       (27'h01F024C),                          // Optimized for IES                                                  
        .PLL1_CFG                       (27'h01F024C),                          // Optimized for IES                                                  
        .PLL_CLKOUT_CFG                 (8'd0),                                 // Optimized for IES                                                   
        .PLL0_DMON_CFG                  (1'b0),                                 // Optimized for IES                                                  
        .PLL1_DMON_CFG                  (1'b0),                                 // Optimized for IES                                      
        .PLL0_FBDIV                     (GTP_QPLL_FBDIV),                       // Optimized for IES                                                  
        .PLL1_FBDIV                     (GTP_QPLL_FBDIV),                       // Optimized for IES                                                   
        .PLL0_FBDIV_45                  (5),                                    // Optimized for IES                                                  
        .PLL1_FBDIV_45                  (5),                                    // Optimized for IES                                                  
        .PLL0_INIT_CFG                  (24'h00001E),                           // Optimized for IES                                                  
        .PLL1_INIT_CFG                  (24'h00001E),                           // Optimized for IES                                                   
        .PLL0_LOCK_CFG                  ( 9'h1E8),                              // Optimized for IES    
        .PLL1_LOCK_CFG                  ( 9'h1E8),                              // Optimized for IES                                                                                                                   
        .PLL0_REFCLK_DIV                (1),                                    // Optimized for IES                                                  
        .PLL1_REFCLK_DIV                (1),                                    // Optimized for IES                                                  
                                                                                                                                     
        //---------- MISC ------------------------------------------------------                                                     
        .BIAS_CFG                       (64'h0000000000050001),                 // Optimized for GES                                                 
      //.COMMON_CFG                     (32'd0),                                //                                                                                                   
        .RSVD_ATTR0                     (16'd0),                                //                                                   
        .RSVD_ATTR1                     (16'd0)                                 //                                                   
    
    )
    model_ap2_tst_gtpe2_common_i 
    (
           
        //---------- Clock -----------------------------------------------------                         
        .GTGREFCLK0                     ( 1'd0),                                //                       
        .GTGREFCLK1                     ( 1'd0),                                //                       
        .GTREFCLK0                      (QPLL_GTGREFCLK),                       //                       
        .GTREFCLK1                      ( 1'd0),                                //                       
        .GTEASTREFCLK0                  ( 1'd0),                                //                       
        .GTEASTREFCLK1                  ( 1'd0),                                //                       
        .GTWESTREFCLK0                  ( 1'd0),                                //                       
        .GTWESTREFCLK1                  ( 1'd0),                                //                       
        .PLL0LOCKDETCLK                 (QPLL_QPLLLOCKDETCLK),                  //                       
        .PLL1LOCKDETCLK                 (QPLL_QPLLLOCKDETCLK),                  //                       
        .PLL0LOCKEN                     ( 1'd1),                                //                       
        .PLL1LOCKEN                     ( 1'd1),                                //                       
        .PLL0REFCLKSEL                  ( 3'd1),                                // Optimized for IES                      
        .PLL1REFCLKSEL                  ( 3'd1),                                // Optimized for IES                      
        .PLLRSVD1                       (16'd0),                                // Optimized for IES                    
        .PLLRSVD2                       ( 5'd0),                                // Optimized for IES                  
        
        .PLL0OUTCLK                     (QPLL_QPLLOUTCLK),                      //                       
        .PLL1OUTCLK                     (),                                     //                       
        .PLL0OUTREFCLK                  (QPLL_QPLLOUTREFCLK),                   //                       
        .PLL1OUTREFCLK                  (),                                     //                       
        .PLL0LOCK                       (QPLL_QPLLLOCK),                        //                       
        .PLL1LOCK                       (),                                     //                       
        .PLL0FBCLKLOST                  (),                                     //                       
        .PLL1FBCLKLOST                  (),                                     //                       
        .PLL0REFCLKLOST                 (),                                     //                       
        .PLL1REFCLKLOST                 (),                                     //                       
        .DMONITOROUT                    (),                                     // 
                                                                                                         
        //---------- Reset -----------------------------------------------------                         
        .PLL0PD                         (cpllpd | QPLL_QPLLPD),                 //                       
        .PLL1PD                         ( 1'd1),                                //                       
        .PLL0RESET                      (cpllrst | QPLL_QPLLRESET),             //                       
        .PLL1RESET                      ( 1'd1),                                //                       
                                                                                                   
        //---------- DRP -------------------------------------------------------                         
        .DRPCLK                         (QPLL_DRPCLK),                          //                       
        .DRPADDR                        (QPLL_DRPADDR),                         //                       
        .DRPEN                          (QPLL_DRPEN),                           //                       
        .DRPDI                          (QPLL_DRPDI),                           //                       
        .DRPWE                          (QPLL_DRPWE),                           //                       
                                                                                                         
        .DRPDO                          (QPLL_DRPDO),                           //                       
        .DRPRDY                         (QPLL_DRPRDY),                          //                       
                                                                                                         
        //---------- Band Gap --------------------------------------------------                         
        .BGBYPASSB                      ( 1'd1),                                // Optimized for IES                      
        .BGMONITORENB                   ( 1'd1),                                // Optimized for IES                      
        .BGPDB                          ( 1'd1),                                // Optimized for IES
        .BGRCALOVRD                     ( 5'd31),                               // Optimized for IES
        .BGRCALOVRDENB                  ( 1'd1),                                // Optimized for IES
        
        //---------- MISC ------------------------------------------------------
        .PMARSVD                        ( 8'd0),                                //
        .RCALENB                        ( 1'd1),                                // Optimized for IES
                                                                               
        .REFCLKOUTMONITOR0              (),                                     //
        .REFCLKOUTMONITOR1              (),                                     //
        .PMARSVDOUT                     ()                                      //  
    
    );
   
    end

else if (PCIE_GT_DEVICE == "GTH") 
    
    //---------- GTH Common ----------------------------------------------------
    begin : gth_common
    
    //---------- GTX Common Module ---------------------------------------------
    GTHE2_COMMON #
    (
       
        //---------- Simulation Attributes -------------------------------------
        .SIM_QPLLREFCLK_SEL             (3'b001),                               //
        .SIM_RESET_SPEEDUP              (PCIE_SIM_MODE),                        //
        .SIM_VERSION                    ("2.0"),                                // 
        
        //---------- Clock Attributes ------------------------------------------
        .QPLL_CFG                       (27'h04801C7),                          // QPLL for Gen3, optimized for GES
        .QPLL_CLKOUT_CFG                ( 4'b1111),                             // Optimized for GES
        .QPLL_COARSE_FREQ_OVRD          ( 6'b010000),                           // 
        .QPLL_COARSE_FREQ_OVRD_EN       ( 1'd0),                                // 
        .QPLL_CP                        (10'h0FF),                              // * Optimized for IES and PCIe PLL BW 
        .QPLL_CP_MONITOR_EN             ( 1'd0),                                //
        .QPLL_DMONITOR_SEL              ( 1'd0),                                //
        .QPLL_FBDIV                     (QPLL_FBDIV),                           // 
        .QPLL_FBDIV_MONITOR_EN          ( 1'd0),                                //
        .QPLL_FBDIV_RATIO               ( 1'd1),                                // Optimized
        .QPLL_INIT_CFG	                (24'h000006),                           // 
        .QPLL_LOCK_CFG                  (16'h05E8),                             // Optimized for IES
        .QPLL_LPF                       ( 4'hD),                                // Optimized for IES, [1:0] = 2'b00 (13.3 KOhm), [1:0] = 2'b01 (57.0 KOhm)
        .QPLL_REFCLK_DIV	              ( 1),                                   // 
        .QPLL_RP_COMP                   ( 1'd0),                                // GTH new
        .QPLL_VTRL_RESET                ( 2'd0),                                // GTH new
    
        //---------- MISC ------------------------------------------------------
        .BIAS_CFG	                      (64'h0000040000001050),                 // Optimized for GES
        .COMMON_CFG	                    (32'd0),                                // 
        .RCAL_CFG                       ( 2'b00),                               // GTH new
        .RSVD_ATTR0                     (16'd0),                                // GTH
        .RSVD_ATTR1                     (16'd0)                                 // GTH    
    )
    model_ap2_tst_gthe2_common_i 
    (
           
        //---------- Clock -----------------------------------------------------
        .GTGREFCLK                      ( 1'd0),                                //    
        .GTREFCLK0                      (QPLL_GTGREFCLK),                       //
        .GTREFCLK1                      ( 1'd0),                                //
        .GTNORTHREFCLK0                 ( 1'd0),                                //
        .GTNORTHREFCLK1                 ( 1'd0),                                //
        .GTSOUTHREFCLK0                 ( 1'd0),                                //
        .GTSOUTHREFCLK1                 ( 1'd0),                                //
        .QPLLLOCKDETCLK                 (QPLL_QPLLLOCKDETCLK),                  //
        .QPLLLOCKEN                     ( 1'd1),                                //
        .QPLLREFCLKSEL                  ( 3'd1),                                //
        .QPLLRSVD1                      (16'd0),                                //
        .QPLLRSVD2                      ( 5'b11111),                            //
                                                                               
        .QPLLOUTCLK                     (QPLL_QPLLOUTCLK),                      //
        .QPLLOUTREFCLK                  (QPLL_QPLLOUTREFCLK),                   //
        .QPLLLOCK                       (QPLL_QPLLLOCK),                        //
        .QPLLFBCLKLOST                  (),                                     //
        .QPLLREFCLKLOST                 (),                                     //
        .QPLLDMONITOR                   (),                                     //
        
        //---------- Reset -----------------------------------------------------
        .QPLLPD                         (QPLL_QPLLPD),                          // 
        .QPLLRESET                      (QPLL_QPLLRESET),                       //
        .QPLLOUTRESET                   ( 1'd0),                                //
        
        //---------- DRP -------------------------------------------------------
        .DRPCLK                         (QPLL_DRPCLK),                          //
        .DRPADDR                        (QPLL_DRPADDR),                         //
        .DRPEN                          (QPLL_DRPEN),                           //
        .DRPDI                          (QPLL_DRPDI),                           //
        .DRPWE                          (QPLL_DRPWE),                           //
                                                                              
        .DRPDO                          (QPLL_DRPDO),                           //
        .DRPRDY                         (QPLL_DRPRDY),                          //
                
        //---------- Band Gap --------------------------------------------------    
        .BGBYPASSB                      ( 1'd1),                                // Optimized for IES
        .BGMONITORENB                   ( 1'd1),                                // Optimized for IES
        .BGPDB                          ( 1'd1),                                // Optimized for IES
        .BGRCALOVRD                     ( 5'd31),                               // Optimized for IES
        .BGRCALOVRDENB                  ( 1'd1),                                // GTH, Optimized for IES
        
        //---------- MISC ------------------------------------------------------
        .PMARSVD                        ( 8'd0),                                //
        .RCALENB                        ( 1'd1),                                // Optimized for IES
                                                                              
        .REFCLKOUTMONITOR               (),                                     //
        .PMARSVDOUT                     ()                                      // GTH
    
    );

    end    
    
else

    //---------- GTX Common ----------------------------------------------------
    begin : gtx_common

    //---------- GTX Common Module ---------------------------------------------
    GTXE2_COMMON #
    (
       
        //---------- Simulation Attributes ------------------------------------- 
        .SIM_QPLLREFCLK_SEL             ( 3'b001),                              //
        .SIM_RESET_SPEEDUP              (PCIE_SIM_MODE),                        //
        .SIM_VERSION                    (PCIE_USE_MODE),                        // 
        
        //---------- Clock Attributes ------------------------------------------
        .QPLL_CFG                       (27'h06801C1),                          // QPLL for Gen3, Optimized for silicon, 
      //.QPLL_CLKOUT_CFG                ( 4'd0),                                //
        .QPLL_COARSE_FREQ_OVRD          ( 6'b010000),                           // 
        .QPLL_COARSE_FREQ_OVRD_EN       ( 1'd0),                                // 
        .QPLL_CP                        (10'h01F),                              // Optimized for Gen3 compliance (Gen1/Gen2 = 10'h1FF) 
        .QPLL_CP_MONITOR_EN             ( 1'd0),                                //
        .QPLL_DMONITOR_SEL              ( 1'd0),                                //
        .QPLL_FBDIV                     (QPLL_FBDIV),                           // 
        .QPLL_FBDIV_MONITOR_EN          ( 1'd0),                                //
        .QPLL_FBDIV_RATIO               ( 1'd1),                                // Optimized for silicon
      //.QPLL_INIT_CFG	                (24'h000006),                           // 
        .QPLL_LOCK_CFG                  (16'h21E8),                             // Optimized for silicon, IES = 16'h01D0, GES 16'h21D0
        .QPLL_LPF                       ( 4'hD),                                // Optimized for silicon, [1:0] = 2'b00 (13.3 KOhm), [1:0] = 2'b01 (57.0 KOhm)
        .QPLL_REFCLK_DIV	              (1),                                    // 
    
        //---------- MISC ------------------------------------------------------
        .BIAS_CFG                       (BIAS_CFG)                              // Optimized for silicon
      //.COMMON_CFG                     (32'd0)                                 //
    
    )
    model_ap2_tst_gtxe2_common_i 
    (
           
        //---------- Clock -----------------------------------------------------
        .GTGREFCLK                      ( 1'd0),                                //
        .GTREFCLK0                      (QPLL_GTGREFCLK),                       //
        .GTREFCLK1                      ( 1'd0),                                //
        .GTNORTHREFCLK0                 ( 1'd0),                                //
        .GTNORTHREFCLK1                 ( 1'd0),                                //
        .GTSOUTHREFCLK0                 ( 1'd0),                                //
        .GTSOUTHREFCLK1                 ( 1'd0),                                //
        .QPLLLOCKDETCLK                 (QPLL_QPLLLOCKDETCLK),                  //
        .QPLLLOCKEN                     ( 1'd1),                                //
        .QPLLREFCLKSEL                  ( 3'd1),                                //
        .QPLLRSVD1                      (16'd0),                                //
        .QPLLRSVD2                      ( 5'b11111),                            //
                                                                               
        .QPLLOUTCLK                     (QPLL_QPLLOUTCLK),                      //
        .QPLLOUTREFCLK                  (QPLL_QPLLOUTREFCLK),                   //
        .QPLLLOCK                       (QPLL_QPLLLOCK),                        //
        .QPLLFBCLKLOST                  (),                                     //
        .QPLLREFCLKLOST                 (),                                     //
        .QPLLDMONITOR                   (),                                     //
        
        //---------- Reset -----------------------------------------------------
        .QPLLPD                         (QPLL_QPLLPD),                          // 
        .QPLLRESET                      (QPLL_QPLLRESET),                       //
        .QPLLOUTRESET                   ( 1'd0),                                //
        
        //---------- DRP -------------------------------------------------------
        .DRPCLK                         (QPLL_DRPCLK),                          //
        .DRPADDR                        (QPLL_DRPADDR),                         //
        .DRPEN                          (QPLL_DRPEN),                           //
        .DRPDI                          (QPLL_DRPDI),                           //
        .DRPWE                          (QPLL_DRPWE),                           //
                                                                               
        .DRPDO                          (QPLL_DRPDO),                           //
        .DRPRDY                         (QPLL_DRPRDY),                          //
                
        //---------- Band Gap --------------------------------------------------    
        .BGBYPASSB                      ( 1'd1),                                //
        .BGMONITORENB                   ( 1'd1),                                //
        .BGPDB                          ( 1'd1),                                //
        .BGRCALOVRD                     ( 5'd31),                               //
        
        //---------- MISC ------------------------------------------------------
        .PMARSVD                        ( 8'd0),                                //
        .RCALENB                        ( 1'd1),                                // Optimized for GES
                                                                               
        .REFCLKOUTMONITOR               ()                                      //
    
    );
    
    end
            
endgenerate

model_ap2_tst_gtp_cpllpd_ovrd model_ap2_tst_cpllPDInst (                                                                                   
        .i_ibufds_gte2(QPLL_CPLLPDREFCLK),                                                                                 
        .o_cpllpd_ovrd(cpllpd),                                                                                       
        .o_cpllreset_ovrd(cpllrst));                       


endmodule

                                              



`timescale 1ns/1ps
module model_ap2_tst_gtp_cpllpd_ovrd (                                                                                        
    input   i_ibufds_gte2,                                                                                     
    output  o_cpllpd_ovrd,                                                                                     
    output  o_cpllreset_ovrd                                                                                   
    );                                                                                                         
    (* equivalent_register_removal="no" *)  reg [95:0] cpllpd_wait = 96'hFFFFFFFFFFFFFFFFFFFFFFFF;             
    (* equivalent_register_removal="no" *)  reg [127:0] cpllreset_wait = 128'h000000000000000000000000000000FF;
    always @(posedge i_ibufds_gte2)                                                                            
    begin                                                                                                      
        cpllpd_wait <= {cpllpd_wait[94:0], 1'b0};                                                              
        cpllreset_wait <= {cpllreset_wait[126:0], 1'b0};                                                       
    end                                                                                                        
    assign o_cpllpd_ovrd = cpllpd_wait[95];                                                                    
    assign o_cpllreset_ovrd = cpllreset_wait[127];                                                             
endmodule



module model_ap2_tst_gt_wrapper #
(
    parameter PCIE_SIM_MODE                 = "FALSE",      // PCIe sim mode
    parameter PCIE_SIM_SPEEDUP              = "FALSE",      // PCIe sim speedup
    parameter PCIE_SIM_TX_EIDLE_DRIVE_LEVEL = "1",          // PCIe sim TX electrical idle drive level
    parameter PCIE_GT_DEVICE                = "GTX",        // PCIe GT device
    parameter PCIE_USE_MODE                 = "3.0",        // PCIe use mode
    parameter PCIE_PLL_SEL                  = "CPLL",       // PCIe PLL select for Gen1/Gen2
    parameter PCIE_LPM_DFE                  = "LPM",        // PCIe LPM or DFE mode for Gen1/Gen2 only
    parameter PCIE_LPM_DFE_GEN3             = "DFE",        // PCIe LPM or DFE mode for Gen3      only
    parameter PCIE_ASYNC_EN                 = "FALSE",      // PCIe async enable
    parameter PCIE_TXBUF_EN                 = "FALSE",      // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_TXSYNC_MODE              = 0,            // PCIe TX sync mode
    parameter PCIE_RXSYNC_MODE              = 0,            // PCIe RX sync mode
    parameter PCIE_CHAN_BOND                = 0,            // PCIe channel bonding mode
    parameter PCIE_CHAN_BOND_EN             = "TRUE",       // PCIe channel bonding enable for Gen1/Gen2 only
    parameter PCIE_LANE                     = 1,            // PCIe number of lane
    parameter PCIE_REFCLK_FREQ              = 0,            // PCIe reference clock frequency
    parameter PCIE_TX_EIDLE_ASSERT_DELAY    = 3'd4,         // PCIe TX electrical idle assert delay
    parameter PCIE_OOBCLK_MODE              = 1,            // PCIe OOB clock mode
    parameter TX_MARGIN_FULL_0              = 7'b1001111,   // 1000 mV
    parameter TX_MARGIN_FULL_1              = 7'b1001110,   // 950 mV
    parameter TX_MARGIN_FULL_2              = 7'b1001101,   // 900 mV
    parameter TX_MARGIN_FULL_3              = 7'b1001100,   // 850 mV
    parameter TX_MARGIN_FULL_4              = 7'b1000011,   // 400 mV
    parameter TX_MARGIN_LOW_0               = 7'b1000101,   // 500 mV
    parameter TX_MARGIN_LOW_1               = 7'b1000110 ,  // 450 mV
    parameter TX_MARGIN_LOW_2               = 7'b1000011,   // 400 mV
    parameter TX_MARGIN_LOW_3               = 7'b1000010 ,  // 350 mV
    parameter TX_MARGIN_LOW_4               = 7'b1000000 ,
    parameter PCIE_DEBUG_MODE               = 0             // PCIe debug mode
)

(    
    //---------- GT User Ports -----------------------------
    input               GT_MASTER,
    input               GT_GEN3, 
    input               GT_RX_CONVERGE,
    
    //---------- GT Clock Ports ----------------------------
    input               GT_GTREFCLK0,
    input               GT_QPLLCLK,
    input               GT_QPLLREFCLK,
    input               GT_TXUSRCLK,
    input               GT_RXUSRCLK,
    input               GT_TXUSRCLK2,
    input               GT_RXUSRCLK2, 
    input               GT_OOBCLK,
    input       [ 1:0]  GT_TXSYSCLKSEL,
    input       [ 1:0]  GT_RXSYSCLKSEL,                
    input               GT_CPLLPDREFCLK,                   
    output              GT_TXOUTCLK,
    output              GT_RXOUTCLK,
    output              GT_CPLLLOCK,
    output              GT_RXCDRLOCK,
    
    //---------- GT Reset Ports ----------------------------
    input               GT_CPLLPD,
    input               GT_CPLLRESET,
    input               GT_TXUSERRDY,
    input               GT_RXUSERRDY,
    input               GT_RESETOVRD,
    input               GT_GTTXRESET,
    input               GT_GTRXRESET,
    input               GT_TXPMARESET,
    input               GT_RXPMARESET,
    input               GT_RXCDRRESET,
    input               GT_RXCDRFREQRESET,
    input               GT_RXDFELPMRESET,
    input               GT_EYESCANRESET,
    input               GT_TXPCSRESET,
    input               GT_RXPCSRESET,
    input               GT_RXBUFRESET,
    
    output              GT_EYESCANDATAERROR,
    output              GT_TXRESETDONE,
    output              GT_RXRESETDONE,
    output              GT_RXPMARESETDONE,
    
    //---------- GT TX Data Ports --------------------------
    input       [31:0]  GT_TXDATA,
    input       [ 3:0]  GT_TXDATAK,
    
    output              GT_TXP,
    output              GT_TXN,
    
    //---------- GT RX Data Ports --------------------------
    input               GT_RXN,
    input               GT_RXP,
    
    output      [31:0]  GT_RXDATA,
    output      [ 3:0]  GT_RXDATAK,
    
    //---------- GT Command Ports --------------------------
    input               GT_TXDETECTRX,
    input               GT_TXELECIDLE,
    input               GT_TXCOMPLIANCE,
    input               GT_RXPOLARITY,
    input       [ 1:0]  GT_TXPOWERDOWN,
    input       [ 1:0]  GT_RXPOWERDOWN,
    input       [ 2:0]  GT_TXRATE,
    input       [ 2:0]  GT_RXRATE,
      
    //---------- GT Electrical Command Ports ---------------
    input       [ 2:0]  GT_TXMARGIN,
    input               GT_TXSWING,
    input               GT_TXDEEMPH,
    input       [ 4:0]  GT_TXPRECURSOR,
    input       [ 6:0]  GT_TXMAINCURSOR,
    input       [ 4:0]  GT_TXPOSTCURSOR,
       
    //---------- GT Status Ports ---------------------------
    output              GT_RXVALID,
    output              GT_PHYSTATUS,
    output              GT_RXELECIDLE,
    output      [ 2:0]  GT_RXSTATUS,
    output      [ 2:0]  GT_RXBUFSTATUS,
    output              GT_TXRATEDONE,
    output              GT_RXRATEDONE,

    output      [7:0]   GT_RXDISPERR,  
    output      [7:0]   GT_RXNOTINTABLE,

    //---------- GT DRP Ports ------------------------------
    input               GT_DRPCLK,
    input       [ 8:0]  GT_DRPADDR,
    input               GT_DRPEN,
    input       [15:0]  GT_DRPDI,
    input               GT_DRPWE,
    
    output      [15:0]  GT_DRPDO,
    output              GT_DRPRDY,
    
    //---------- GT TX Sync Ports --------------------------
    input               GT_TXPHALIGN,     
    input               GT_TXPHALIGNEN,  
    input               GT_TXPHINIT, 
    input               GT_TXDLYBYPASS,
    input               GT_TXDLYSRESET,
    input               GT_TXDLYEN,       
    
    output              GT_TXDLYSRESETDONE,
    output              GT_TXPHINITDONE,  
    output              GT_TXPHALIGNDONE,
    
    input               GT_TXPHDLYRESET,
    input               GT_TXSYNCMODE,                      // GTH
    input               GT_TXSYNCIN,                        // GTH
    input               GT_TXSYNCALLIN,                     // GTH
        
    output              GT_TXSYNCOUT,                       // GTH                                                                        
    output              GT_TXSYNCDONE,                      // GTH                                                                        
                                                                            
    //---------- GT RX Sync Ports --------------------------
    input               GT_RXPHALIGN,
    input               GT_RXPHALIGNEN,
    input               GT_RXDLYBYPASS,
    input               GT_RXDLYSRESET,
    input               GT_RXDLYEN,
    input               GT_RXDDIEN,
    
    output              GT_RXDLYSRESETDONE,
    output              GT_RXPHALIGNDONE,    
    
    input               GT_RXSYNCMODE,                      // GTH
    input               GT_RXSYNCIN,                        // GTH
    input               GT_RXSYNCALLIN,                     // GTH
    
    output              GT_RXSYNCOUT,                       // GTH
    output              GT_RXSYNCDONE,                      // GTH
    
    //---------- GT Comma Alignment Ports ------------------
    input               GT_RXSLIDE,
    
    output              GT_RXCOMMADET,                        
    output      [ 3:0]  GT_RXCHARISCOMMA,                      
    output              GT_RXBYTEISALIGNED,                   
    output              GT_RXBYTEREALIGN,                     
    
    //---------- GT Channel Bonding Ports ------------------
    input               GT_RXCHBONDEN,
    input       [ 4:0]  GT_RXCHBONDI,
    input       [ 2:0]  GT_RXCHBONDLEVEL,
    input               GT_RXCHBONDMASTER,
    input               GT_RXCHBONDSLAVE,
    
    output              GT_RXCHANISALIGNED,
    output      [ 4:0]  GT_RXCHBONDO,
    
    //---------- GT PRBS/Loopback Ports --------------------
    input       [ 2:0]  GT_TXPRBSSEL,
    input       [ 2:0]  GT_RXPRBSSEL,
    input               GT_TXPRBSFORCEERR,
    input               GT_RXPRBSCNTRESET,
    input       [ 2:0]  GT_LOOPBACK,
    
    output              GT_RXPRBSERR,
    
    //---------- GT Debug Ports ----------------------------
    output      [14:0]  GT_DMONITOROUT

);

    //---------- Internal Signals --------------------------
    wire        [ 2:0]  txoutclksel;
    wire        [ 2:0]  rxoutclksel;
    wire        [63:0]  rxdata;
    wire        [ 7:0]  rxdatak;
    wire        [ 7:0]  rxchariscomma;
    wire rxlpmen;
    wire        [14:0]  dmonitorout;
    wire                dmonitorclk;

    wire cpllpd;
    wire cpllrst;

    //---------- Select CPLL and Clock Dividers ------------
    localparam          CPLL_REFCLK_DIV = 1;
    localparam          CPLL_FBDIV_45   = 5;
    localparam          CPLL_FBDIV      = (PCIE_REFCLK_FREQ == 2) ?  2 : 
                                          (PCIE_REFCLK_FREQ == 1) ?  4 : 5;
    localparam          OUT_DIV         = (PCIE_PLL_SEL == "QPLL") ? 4 : 2;                                                     
    localparam          CLK25_DIV       = (PCIE_REFCLK_FREQ == 2) ? 10 : 
                                          (PCIE_REFCLK_FREQ == 1) ?  5 : 4;
    
    //---------- Select IES vs. GES ------------------------
    localparam          CLKMUX_PD = ((PCIE_USE_MODE == "1.0") || (PCIE_USE_MODE == "1.1")) ?  1'd0      :  1'd1;
    
    //---------- Select GTP CPLL configuration -------------
    //  PLL0/1_CFG[ 5:2] = CP1 : [    8, 4, 2, 1] units
    //  PLL0/1_CFG[10:6] = CP2 : [16, 8, 4, 2, 1] units
    //  CP2/CP1 = 2 to 3  
    //  (8/4=2)    = 27'h01F0210 = 0000_0001_1111_0000_0010_0001_0000
    //  (9/3=3)    = 27'h01F024C = 0000_0001_1111_0000_0010_0100_1100
    //  (8/3=2.67) = 27'h01F020C = 0000_0001_1111_0000_0010_0000_1100
    //  (7/3=2.33) = 27'h01F01CC = 0000_0001_1111_0000_0001_1100_1100
    //  (6/3=2)    = 27'h01F018C = 0000_0001_1111_0000_0001_1000_1100
    //  (5/3=1.67) = 27'h01F014C = 0000_0001_1111_0000_0001_0100_1100
    //  (6/2=3)    = 27'h01F0188 = 0000_0001_1111_0000_0001_1000_1000
    //---------- Select GTX CPLL configuration -------------
    //  CPLL_CFG[ 5: 2]  = CP1 : [    8, 4, 2, 1] units 
    //  CPLL_CFG[22:18]  = CP2 : [16, 8, 4, 2, 1] units
    //  CP2/CP1 = 2 to 3 
    //  (9/3=3)    = 1010_0100_0000_0111_1100_1100
    //------------------------------------------------------
    localparam          CPLL_CFG  = ((PCIE_USE_MODE == "1.0") || (PCIE_USE_MODE == "1.1")) ? 24'hB407CC : 24'hA407CC;
    
    //---------- Select TX XCLK ----------------------------      
    //  TXOUT for TX Buffer Use     
    //  TXUSR for TX Buffer Bypass  
    //------------------------------------------------------                                            
    localparam          TX_XCLK_SEL = (PCIE_TXBUF_EN == "TRUE") ? "TXOUT" : "TXUSR";
                                                   
    //---------- Select TX Receiver Detection Configuration 
    localparam          TX_RXDETECT_CFG = (PCIE_REFCLK_FREQ == 2) ? 14'd250 : 
                                          (PCIE_REFCLK_FREQ == 1) ? 14'd125 : 14'd100;
    localparam          TX_RXDETECT_REF = (((PCIE_USE_MODE == "1.0") || (PCIE_USE_MODE == "1.1")) && (PCIE_SIM_MODE == "FALSE")) ? 3'b000 : 3'b011;                                                                 
                                                      
    //---------- Select PCS_RSVD_ATTR ----------------------
    //  [0]: 1 = enable latch when bypassing TX buffer, 0 = disable latch when using TX buffer 
    //  [1]: 1 = enable manual TX sync,                 0 = enable auto TX sync
    //  [2]: 1 = enable manual RX sync,                 0 = enable auto RX sync
    //  [3]: 1 = select external clock for OOB          0 = select reference clock for OOB    
    //  [6]: 1 = enable DMON                            0 = disable DMON     
    //  [7]: 1 = filter stale TX[P/N] data when exiting TX electrical idle
    //  [8]: 1 = power up OOB                           0 = power down OOB
    //------------------------------------------------------
    localparam          OOBCLK_SEL    = (PCIE_OOBCLK_MODE == 0) ? 1'd0  : 1'd1;      // GTX
    localparam          RXOOB_CLK_CFG = (PCIE_OOBCLK_MODE == 0) ? "PMA" : "FABRIC";  // GTH/GTP
    
    localparam          PCS_RSVD_ATTR = ((PCIE_USE_MODE == "1.0")                           && (PCIE_TXBUF_EN == "FALSE")) ? {44'h0000000001C, OOBCLK_SEL, 3'd1} :
                                        ((PCIE_USE_MODE == "1.0")                           && (PCIE_TXBUF_EN == "TRUE" )) ? {44'h0000000001C, OOBCLK_SEL, 3'd0} : 
                                        ((PCIE_RXSYNC_MODE == 0) && (PCIE_TXSYNC_MODE == 0) && (PCIE_TXBUF_EN == "FALSE")) ? {44'h0000000001C, OOBCLK_SEL, 3'd7} : 
                                        ((PCIE_RXSYNC_MODE == 0) && (PCIE_TXSYNC_MODE == 0) && (PCIE_TXBUF_EN == "TRUE" )) ? {44'h0000000001C, OOBCLK_SEL, 3'd6} :   
                                        ((PCIE_RXSYNC_MODE == 0) && (PCIE_TXSYNC_MODE == 1) && (PCIE_TXBUF_EN == "FALSE")) ? {44'h0000000001C, OOBCLK_SEL, 3'd5} : 
                                        ((PCIE_RXSYNC_MODE == 0) && (PCIE_TXSYNC_MODE == 1) && (PCIE_TXBUF_EN == "TRUE" )) ? {44'h0000000001C, OOBCLK_SEL, 3'd4} : 
                                        ((PCIE_RXSYNC_MODE == 1) && (PCIE_TXSYNC_MODE == 0) && (PCIE_TXBUF_EN == "FALSE")) ? {44'h0000000001C, OOBCLK_SEL, 3'd3} : 
                                        ((PCIE_RXSYNC_MODE == 1) && (PCIE_TXSYNC_MODE == 0) && (PCIE_TXBUF_EN == "TRUE" )) ? {44'h0000000001C, OOBCLK_SEL, 3'd2} : 
                                        ((PCIE_RXSYNC_MODE == 1) && (PCIE_TXSYNC_MODE == 1) && (PCIE_TXBUF_EN == "FALSE")) ? {44'h0000000001C, OOBCLK_SEL, 3'd1} : 
                                        ((PCIE_RXSYNC_MODE == 1) && (PCIE_TXSYNC_MODE == 1) && (PCIE_TXBUF_EN == "TRUE" )) ? {44'h0000000001C, OOBCLK_SEL, 3'd0} : {44'h0000000001C, OOBCLK_SEL, 3'd7};                                      
                             
    //---------- Select RXCDR_CFG --------------------------
    
    //---------- GTX Note ----------------------------------
    // For GTX PCIe Gen1/Gen2 with 8B/10B, the following CDR setting may provide more margin
    // Async 72'h03_8000_23FF_1040_0020
    // Sync: 72'h03_0000_23FF_1040_0020   
    //------------------------------------------------------      
    
    localparam          RXCDR_CFG_GTX = ((PCIE_USE_MODE == "1.0") || (PCIE_USE_MODE == "1.1")) ? 
                                        ((PCIE_ASYNC_EN == "TRUE") ? 72'b0000_0010_0000_0111_1111_1110_0010_0000_0110_0000_0010_0001_0001_0000_0000000000010000
                                                                   : 72'h11_07FE_4060_0104_0000):   // IES setting
                                        ((PCIE_ASYNC_EN == "TRUE") ? 72'h03_8000_23FF_1020_0020     // 
                                                                   : 72'h03_0000_23FF_1020_0020);   // optimized for GES silicon                                                                                
                            
    localparam          RXCDR_CFG_GTH = (PCIE_USE_MODE == "2.0") ? 
                                        ((PCIE_ASYNC_EN == "TRUE") ? 83'h0_0011_07FE_4060_2104_1010   
                                                                   : 83'h0_0011_07FE_4060_0104_1010):  // Optimized for IES silicon
                                        ((PCIE_ASYNC_EN == "TRUE") ? 83'h0_0020_07FE_2000_C208_8018   
                                                                   : 83'h0_0020_07FE_2000_C208_0018);  // Optimized for 1.2 silicon     
                                                                                 
    localparam          RXCDR_CFG_GTP = ((PCIE_ASYNC_EN == "TRUE") ? 83'h0_0001_07FE_4060_2104_1010
                                                                   : 83'h0_0001_07FE_4060_0104_1010);  // Optimized for IES silicon
                   
                         
                                                                                           
                            
    //---------- Select TX and RX Sync Mode ----------------                                            
    localparam          TXSYNC_OVRD      = (PCIE_TXSYNC_MODE == 1) ? 1'd0 : 1'd1;                             
    localparam          RXSYNC_OVRD      = (PCIE_TXSYNC_MODE == 1) ? 1'd0 : 1'd1;     
                                                                          
    localparam          TXSYNC_MULTILANE = (PCIE_LANE == 1) ? 1'd0 : 1'd1;  
    localparam          RXSYNC_MULTILANE = (PCIE_LANE == 1) ? 1'd0 : 1'd1;                                             
                                       
    //---------- Select Clock Correction Min and Max Latency
    //  CLK_COR_MIN_LAT = Larger of (2 * RXCHBONDLEVEL + 13) or (CHAN_BOND_MAX_SKEW + 11)
    //                  = 13 when PCIE_LANE = 1
    //  CLK_COR_MAX_LAT = CLK_COR_MIN_LAT + CLK_COR_SEQ_LEN + 1
    //                  = CLK_COR_MIN_LAT + 2
    //------------------------------------------------------
   
    //---------- CLK_COR_MIN_LAT Look-up Table -------------
    // Lane | One-Hop  | Daisy-Chain | Binary-Tree
    //------------------------------------------------------
    //    0 |       13 |       13    |       13
    //    1 | 15 to 18 | 15 to 18    | 15 to 18
    //    2 | 15 to 18 | 17 to 18    | 15 to 18
    //    3 | 15 to 18 |       19    | 17 to 18
    //    4 | 15 to 18 |       21    | 17 to 18
    //    5 | 15 to 18 |       23    |       19
    //    6 | 15 to 18 |       25    |       19
    //    7 | 15 to 18 |       27    |       21
    //------------------------------------------------------
    
    localparam          CLK_COR_MIN_LAT = ((PCIE_LANE == 8) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 27 : 21) : 
                                          ((PCIE_LANE == 7) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 25 : 19) : 
                                          ((PCIE_LANE == 6) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 23 : 19) : 
                                          ((PCIE_LANE == 5) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 21 : 18) : 
                                          ((PCIE_LANE == 4) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 19 : 18) :
                                          ((PCIE_LANE == 3) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 18 : 18) :
                                          ((PCIE_LANE == 2) && (PCIE_CHAN_BOND != 0) && (PCIE_CHAN_BOND_EN == "TRUE"))  ? ((PCIE_CHAN_BOND == 1) ? 18 : 18) :
                                          ((PCIE_LANE == 1)                          || (PCIE_CHAN_BOND_EN == "FALSE")) ? 13 : 18; 
                                           
    localparam          CLK_COR_MAX_LAT = CLK_COR_MIN_LAT + 2;                                                     
    
    //---------- Simulation Speedup ------------------------
  //localparam          CFOK_CFG_GTH = (PCIE_SIM_MODE == "TRUE") ? 42'h240_0004_0F80 : 42'h248_0004_0E80;  // [8] : 1 = Skip CFOK
  //localparam          CFOK_CFG_GTP = (PCIE_SIM_MODE == "TRUE") ? 43'h000_0000_0000 : 43'h000_0000_0100;  // [2] : 1 = Skip CFOK

    //---------- Select [TX/RX]OUTCLK ----------------------
    assign txoutclksel = GT_MASTER ? 3'd3 : 3'd0;
    assign rxoutclksel = ((PCIE_DEBUG_MODE == 1) || ((PCIE_ASYNC_EN == "TRUE") && GT_MASTER)) ? 3'd2 : 3'd0;
 
    //---------- Select DFE vs. LPM ------------------------
    //  Gen1/2 = Use LPM by default.  Option to use DFE.
    //  Gen3   = Use DFE by default.  Option to use LPM.
    //------------------------------------------------------
    assign rxlpmen = GT_GEN3 ? ((PCIE_LPM_DFE_GEN3 == "LPM") ? 1'd1 : 1'd0) : ((PCIE_LPM_DFE == "LPM") ? 1'd1 : 1'd0);
    

 
//---------- Generate DMONITOR Clock Buffer for Debug ------  
generate if (PCIE_DEBUG_MODE == 1)
 
    begin : dmonitorclk_i
    //---------- DMONITOR CLK ------------------------------
    BUFG dmonitorclk_i
    (
        //---------- Input ---------------------------------
        .I                              (dmonitorout[7]),   
        //---------- Output --------------------------------
        .O                              (dmonitorclk)
    ); 
    end
    
else

    begin : dmonitorclk_i_disable
    assign dmonitorclk = 1'd0;
    end
    
endgenerate

   
model_ap2_tst_gtx_cpllpd_ovrd cpllPDInst (
   .i_ibufds_gte2(GT_CPLLPDREFCLK),
   .o_cpllpd_ovrd(cpllpd),
   .o_cpllreset_ovrd(cpllrst));
 
//---------- Select GTX or GTH or GTP ------------------------------------------
//  Notes  :  Attributes that are commented out always use the GT default settings
//------------------------------------------------------------------------------
generate if (PCIE_GT_DEVICE == "GTP") 

    begin : gtp_channel

    //---------- GTP Channel Module --------------------------------------------
    GTPE2_CHANNEL #
    (
                
        //---------- Simulation Attributes -------------------------------------
        .SIM_RESET_SPEEDUP              (PCIE_SIM_SPEEDUP),                     //
        .SIM_RECEIVER_DETECT_PASS       ("TRUE"),                               //    
        .SIM_TX_EIDLE_DRIVE_LEVEL       (PCIE_SIM_TX_EIDLE_DRIVE_LEVEL),        // 
        .SIM_VERSION                    (PCIE_USE_MODE),                        //
                                                                                 
        //---------- Clock Attributes ------------------------------------------                                      
        .TXOUT_DIV                      (OUT_DIV),                              //
        .RXOUT_DIV                      (OUT_DIV),                              // 
        .TX_CLK25_DIV                   (CLK25_DIV),                            //
        .RX_CLK25_DIV                   (CLK25_DIV),                            //
      //.TX_CLKMUX_EN                   ( 1'b1),                                // GTP rename
      //.RX_CLKMUX_EN                   ( 1'b1),                                // GTP rename
        .TX_XCLK_SEL                    (TX_XCLK_SEL),                          // TXOUT = use TX buffer, TXUSR = bypass TX buffer
        .RX_XCLK_SEL                    ("RXREC"),                              // RXREC = use RX buffer, RXUSR = bypass RX buffer
      //.OUTREFCLK_SEL_INV              ( 2'b11),                               //
                                                                                 
        //---------- Reset Attributes ------------------------------------------                
        .TXPCSRESET_TIME                ( 5'b00001),                            //
        .RXPCSRESET_TIME                ( 5'b00001),                            //
        .TXPMARESET_TIME                ( 5'b00011),                            //
        .RXPMARESET_TIME                ( 5'b00011),                            // Optimized for sim
      //.RXISCANRESET_TIME              ( 5'b00001),                            //
                                                                                 
        //---------- TX Data Attributes ----------------------------------------                
        .TX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        
        //---------- RX Data Attributes ----------------------------------------                
        .RX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        
        //---------- Command Attributes ----------------------------------------                
        .TX_RXDETECT_CFG                (TX_RXDETECT_CFG),                      // 
        .TX_RXDETECT_REF                ( 3'b011),                              // 
        .RX_CM_SEL                      ( 2'd3),                                // 0 = AVTT, 1 = GND, 2 = Float, 3 = Programmable
        .RX_CM_TRIM	                    ( 4'b1010),                             // Select 800mV, Changed from 3 to 4-bits, optimized for IES
        .TX_EIDLE_ASSERT_DELAY          (PCIE_TX_EIDLE_ASSERT_DELAY),           // Optimized for sim
        .TX_EIDLE_DEASSERT_DELAY        ( 3'b010),                              // Optimized for sim
      //.PD_TRANS_TIME_FROM_P2          (12'h03C),                              //
        .PD_TRANS_TIME_NONE_P2          ( 8'h09),                               //
      //.PD_TRANS_TIME_TO_P2            ( 8'h64),                               //
      //.TRANS_TIME_RATE                ( 8'h0E),                               //
                                                                                 
        //---------- Electrical Command Attributes -----------------------------                
        .TX_DRIVE_MODE                  ("PIPE"),                               // Gen1/Gen2 = PIPE, Gen3 = PIPEGEN3
        .TX_DEEMPH0                     ( 5'b10100),                            //  6.0 dB
        .TX_DEEMPH1                     ( 5'b01011),                            //  3.5 dB
        .TX_MARGIN_FULL_0               ( 7'b1001111),                          // 1000 mV
        .TX_MARGIN_FULL_1               ( 7'b1001110),                          //  950 mV
        .TX_MARGIN_FULL_2               ( 7'b1001101),                          //  900 mV
        .TX_MARGIN_FULL_3               ( 7'b1001100),                          //  850 mV
        .TX_MARGIN_FULL_4               ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_0                ( 7'b1000101),                          //  500 mV
        .TX_MARGIN_LOW_1                ( 7'b1000110),                          //  450 mV
        .TX_MARGIN_LOW_2                ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_3                ( 7'b1000010),                          //  350 mV
        .TX_MARGIN_LOW_4                ( 7'b1000000),                          //  250 mV
        .TX_MAINCURSOR_SEL              ( 1'b0),                                //
        .TX_PREDRIVER_MODE              ( 1'b0),                                // GTP
                                                                                
        //---------- Status Attributes -----------------------------------------                
      //.RX_SIG_VALID_DLY               ( 4),                                   // CHECK
                                                                                 
        //---------- DRP Attributes --------------------------------------------                
                          
        //---------- PCS Attributes --------------------------------------------                
        .PCS_PCIE_EN                    ("TRUE"),                               // PCIe
        .PCS_RSVD_ATTR                  (48'h0000_0000_0100),                   // [8] : 1 = OOB power-up
                                                                                 
         //---------- PMA Attributes ------------------------------------------- 
      //.CLK_COMMON_SWING               ( 1'b0),                                // GTP new              
      //.PMA_RSV                        (32'd0),                                // 
        .PMA_RSV2                       (32'h00002040),                         // Optimized for GES
      //.PMA_RSV3                       ( 2'd0),                                // 
      //.PMA_RSV4                       ( 4'd0),                                // Changed from 15 to 4-bits
      //.PMA_RSV5                       ( 1'd0),                                // Changed from 4 to 1-bit
      //.PMA_RSV6                       ( 1'd0),                                // GTP new
      //.PMA_RSV7                       ( 1'd0),                                // GTP new
        .RX_BIAS_CFG                    (16'h0F33),                             // Optimized for IES
        .TERM_RCAL_CFG                  (15'b100001000010000),                  // Optimized for IES
        .TERM_RCAL_OVRD                 ( 3'b000),                              // Optimized for IES 
                                             
         //---------- TX PI ----------------------------------------------------                                              
      //.TXPI_CFG0                      ( 2'd0),                                //                                            
      //.TXPI_CFG1                      ( 2'd0),                                //                                            
      //.TXPI_CFG2                      ( 2'd0),                                //                                            
      //.TXPI_CFG3                      ( 1'd0),                                //                                            
      //.TXPI_CFG4                      ( 1'd0),                                //                                            
      //.TXPI_CFG5                      ( 3'd000),                              //                                            
      //.TXPI_GREY_SEL                  ( 1'd0),                                //                                            
      //.TXPI_INVSTROBE_SEL             ( 1'd0),                                //                                            
      //.TXPI_PPMCLK_SEL                ("TXUSRCLK2"),                          //                                            
      //.TXPI_PPM_CFG                   ( 8'd0),                                //                                            
      //.TXPI_SYNFREQ_PPM               ( 3'd0),                                //                                            
                                                                                                                               
        //---------- RX PI -----------------------------------------------------                                              
        .RXPI_CFG0                      ( 3'd0),                                // Changed from 3 to 2-bits, Optimized for IES                                           
        .RXPI_CFG1                      ( 1'd1),                                // Changed from 2 to 1-bits, Optimized for IES                                          
        .RXPI_CFG2                      ( 1'd1),                                // Changed from 2 to 1-bits, Optimized for IES                                                      
                                             
       //---------- CDR Attributes ---------------------------------------------
      //.RXCDR_CFG                      (72'b0000_001000000_11111_11111_001000000_011_0000111_000_001000_010000_100000000000000),  // CHECK  
        .RXCDR_CFG                      (RXCDR_CFG_GTP),       // Optimized for IES                       
        .RXCDR_LOCK_CFG                 ( 6'b010101),                           // [5:3] Window Refresh, [2:1] Window Size, [0] Enable Detection (sensitive lock = 6'b111001)  CHECK
        .RXCDR_HOLD_DURING_EIDLE        ( 1'd1),                                // Hold  RX CDR           on electrical idle for Gen1/Gen2
        .RXCDR_FR_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR frequency on electrical idle for Gen3
        .RXCDR_PH_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR phase     on electrical idle for Gen3
      //.RXCDRFREQRESET_TIME            ( 5'b00001),                            // 
      //.RXCDRPHRESET_TIME              ( 5'b00001),                            // 
                                  
        //---------- LPM Attributes --------------------------------------------               
      //.RXLPMRESET_TIME                ( 7'b0001111),                          // GTP new
      //.RXLPM_BIAS_STARTUP_DISABLE     ( 1'b0),                                // GTP new
        .RXLPM_CFG                      ( 4'b0110),                             // GTP new, optimized for IES
      //.RXLPM_CFG1                     ( 1'b0),                                // GTP new
      //.RXLPM_CM_CFG                   ( 1'b0),                                // GTP new
        .RXLPM_GC_CFG                   ( 9'b111100010),                        // GTP new, optimized for IES
        .RXLPM_GC_CFG2                  ( 3'b001),                              // GTP new, optimized for IES
      //.RXLPM_HF_CFG                   (14'b00001111110000),                   //
        .RXLPM_HF_CFG2                  ( 5'b01010),                            // GTP new
      //.RXLPM_HF_CFG3                  ( 4'b0000),                             // GTP new
        .RXLPM_HOLD_DURING_EIDLE        ( 1'b1),                                // GTP new
        .RXLPM_INCM_CFG                 ( 1'b1),                                // GTP new, optimized for IES
        .RXLPM_IPCM_CFG                 ( 1'b0),                                // GTP new, optimized for IES
      //.RXLPM_LF_CFG                   (18'b000000001111110000),               // 
        .RXLPM_LF_CFG2                  ( 5'b01010),                            // GTP new, optimized for IES
        .RXLPM_OSINT_CFG                ( 3'b100),                              // GTP new, optimized for IES
                                                                           
        //---------- OS Attributes ---------------------------------------------
        .RX_OS_CFG                      (13'h0080),                             // CHECK
        .RXOSCALRESET_TIME              (5'b00011),                             // Optimized for IES
        .RXOSCALRESET_TIMEOUT           (5'b00000),                             // Disable timeout, Optimized for IES     
                                                                                 
        //---------- Eye Scan Attributes --------------------------------------- 
      //.ES_CLK_PHASE_SEL               ( 1'b0),                                //
      //.ES_CONTROL                     ( 6'd0),                                //
      //.ES_ERRDET_EN                   ("FALSE"),                              //
        .ES_EYE_SCAN_EN                 ("FALSE"),                               // 
      //.ES_HORZ_OFFSET                 (12'd0),                                //
      //.ES_PMA_CFG                     (10'd0),                                //
      //.ES_PRESCALE                    ( 5'd0),                                //
      //.ES_QUAL_MASK                   (80'd0),                                //
      //.ES_QUALIFIER                   (80'd0),                                //
      //.ES_SDATA_MASK                  (80'd0),                                //
      //.ES_VERT_OFFSET                 ( 9'd0),                                //
                                                                                 
        //---------- TX Buffer Attributes --------------------------------------               
        .TXBUF_EN                       (PCIE_TXBUF_EN),                        // 
        .TXBUF_RESET_ON_RATE_CHANGE     ("TRUE"),                               //
                                                                                 
        //---------- RX Buffer Attributes --------------------------------------                
        .RXBUF_EN                       ("TRUE"),                               //
      //.RX_BUFFER_CFG                  ( 6'd0),                                //
        .RX_DEFER_RESET_BUF_EN          ("TRUE"),                               // 
        .RXBUF_ADDR_MODE                ("FULL"),                               //
        .RXBUF_EIDLE_HI_CNT	            ( 4'd4),                                // Optimized for sim
        .RXBUF_EIDLE_LO_CNT	            ( 4'd0),                                // Optimized for sim
        .RXBUF_RESET_ON_CB_CHANGE       ("TRUE"),                               //
        .RXBUF_RESET_ON_COMMAALIGN      ("FALSE"),                              //
        .RXBUF_RESET_ON_EIDLE           ("TRUE"),                               // PCIe
        .RXBUF_RESET_ON_RATE_CHANGE     ("TRUE"),                               //
        .RXBUF_THRESH_OVRD              ("FALSE"),                              //
        .RXBUF_THRESH_OVFLW             (61),                                   //
        .RXBUF_THRESH_UNDFLW            ( 4),                                   //
      //.RXBUFRESET_TIME                ( 5'b00001),                            //
                                                                                 
        //---------- TX Sync Attributes ----------------------------------------                
        .TXPH_CFG                       (16'h0780),                             // 
        .TXPH_MONITOR_SEL               ( 5'd0),                                // 
        .TXPHDLY_CFG                    (24'h084020),                           // [19] : 1 = full range, 0 = half range
        .TXDLY_CFG                      (16'h001F),                             // 
        .TXDLY_LCFG	                    ( 9'h030),                              // 
        .TXDLY_TAP_CFG                  (16'd0),                                // 
                 
        .TXSYNC_OVRD                    (TXSYNC_OVRD),                          //
        .TXSYNC_MULTILANE               (TXSYNC_MULTILANE),                     //
        .TXSYNC_SKIP_DA                 (1'b0),                                 //
                                                                                 
        //---------- RX Sync Attributes ----------------------------------------            
        .RXPH_CFG                       (24'd0),                                //
        .RXPH_MONITOR_SEL               ( 5'd0),                                //
        .RXPHDLY_CFG                    (24'h004020),                           // [19] : 1 = full range, 0 = half range
        .RXDLY_CFG                      (16'h001F),                             // 
        .RXDLY_LCFG	                    ( 9'h030),                              //
        .RXDLY_TAP_CFG                  (16'd0),                                //
        .RX_DDI_SEL	                    ( 6'd0),                                //
            
        .RXSYNC_OVRD                    (RXSYNC_OVRD),                          //    
        .RXSYNC_MULTILANE               (RXSYNC_MULTILANE),                     //
        .RXSYNC_SKIP_DA                 (1'b0),                                 //
                                                                                 
        //---------- Comma Alignment Attributes --------------------------------            
        .ALIGN_COMMA_DOUBLE             ("FALSE"),                              //   
        .ALIGN_COMMA_ENABLE             (10'b1111111111),                       // PCIe
        .ALIGN_COMMA_WORD               ( 1),                                   //
        .ALIGN_MCOMMA_DET               ("TRUE"),                               //
        .ALIGN_MCOMMA_VALUE             (10'b1010000011),                       //
        .ALIGN_PCOMMA_DET               ("TRUE"),                               //
        .ALIGN_PCOMMA_VALUE             (10'b0101111100),                       //
        .DEC_MCOMMA_DETECT              ("TRUE"),                               //
        .DEC_PCOMMA_DETECT              ("TRUE"),                               //
        .DEC_VALID_COMMA_ONLY           ("FALSE"),                              // PCIe
        .SHOW_REALIGN_COMMA             ("FALSE"),                              // PCIe
        .RXSLIDE_AUTO_WAIT              ( 7),                                   // 
        .RXSLIDE_MODE                   ("PMA"),                                // PCIe
                                                                                 
        //---------- Channel Bonding Attributes --------------------------------                
        .CHAN_BOND_KEEP_ALIGN           ("TRUE"),                               // PCIe
        .CHAN_BOND_MAX_SKEW             ( 7),                                   // 
        .CHAN_BOND_SEQ_LEN              ( 4),                                   // PCIe
        .CHAN_BOND_SEQ_1_ENABLE         ( 4'b1111),                             //
        .CHAN_BOND_SEQ_1_1              (10'b0001001010),                       // D10.2 (4A) - TS1 
        .CHAN_BOND_SEQ_1_2              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_3              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .CHAN_BOND_SEQ_2_USE            ("TRUE"),                               // PCIe
        .CHAN_BOND_SEQ_2_ENABLE         (4'b1111),                              //
        .CHAN_BOND_SEQ_2_1              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_2              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_3              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .FTS_DESKEW_SEQ_ENABLE          ( 4'b1111),                             // 
        .FTS_LANE_DESKEW_EN             ("TRUE"),                               // PCIe
        .FTS_LANE_DESKEW_CFG            ( 4'b1111),                             // 
                                                                                 
        //---------- Clock Correction Attributes -------------------------------        
        .CBCC_DATA_SOURCE_SEL           ("DECODED"),                            //
        .CLK_CORRECT_USE                ("TRUE"),                               //
        .CLK_COR_KEEP_IDLE              ("TRUE"),                               // PCIe
        .CLK_COR_MAX_LAT                (CLK_COR_MAX_LAT),                      // 
        .CLK_COR_MIN_LAT                (CLK_COR_MIN_LAT),                      // 
        .CLK_COR_PRECEDENCE             ("TRUE"),                               //
        .CLK_COR_REPEAT_WAIT            ( 0),                                   // 
        .CLK_COR_SEQ_LEN                ( 1),                                   //
        .CLK_COR_SEQ_1_ENABLE           ( 4'b1111),                             //
        .CLK_COR_SEQ_1_1                (10'b0100011100),                       // K28.0 (1C) - SKP
        .CLK_COR_SEQ_1_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_4                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_ENABLE           ( 4'b0000),                             // Disabled
        .CLK_COR_SEQ_2_USE              ("FALSE"),                              //
        .CLK_COR_SEQ_2_1                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_4                (10'b0000000000),                       // Disabled
                                                                                 
        //---------- 8b10b Attributes ------------------------------------------                
        .RX_DISPERR_SEQ_MATCH           ("TRUE"),                               //
                                                                                 
        //---------- 64b/66b & 64b/67b Attributes ------------------------------                
        .GEARBOX_MODE                   ( 3'd0),                                //
        .TXGEARBOX_EN                   ("FALSE"),                              //
        .RXGEARBOX_EN                   ("FALSE"),                              //
                                                                                 
       //---------- PRBS & Loopback Attributes ---------------------------------      
        .LOOPBACK_CFG                    ( 1'd0),                               // Enable latch when bypassing TX buffer, equivalent to GTX PCS_RSVD_ATTR[0]      
        .RXPRBS_ERR_LOOPBACK             ( 1'd0),                               //
        .TX_LOOPBACK_DRIVE_HIZ           ("FALSE"),                             //
                                                                                 
       //---------- OOB & SATA Attributes --------------------------------------                
        .TXOOB_CFG                      ( 1'd1),                                // Filter stale TX data when exiting TX electrical idle, equivalent to GTX PCS_RSVD_ATTR[7]
      //.RXOOB_CFG                      ( 7'b0000110),                          //
        .RXOOB_CLK_CFG                  (RXOOB_CLK_CFG),                        // 
      //.SAS_MAX_COM                    (64),                                   //
      //.SAS_MIN_COM                    (36),                                   //
      //.SATA_BURST_SEQ_LEN             ( 4'b1111),                             //
      //.SATA_BURST_VAL                 ( 3'b100),                              //
      //.SATA_PLL_CFG                   ("VCO_3000MHZ"),                        //
      //.SATA_EIDLE_VAL                 ( 3'b100),                              //
      //.SATA_MAX_BURST                 ( 8),                                   //
      //.SATA_MAX_INIT                  (21),                                   //
      //.SATA_MAX_WAKE                  ( 7),                                   //
      //.SATA_MIN_BURST                 ( 4),                                   //
      //.SATA_MIN_INIT                  (12),                                   //
      //.SATA_MIN_WAKE                  ( 4),                                   //  
                                                                                 
        //---------- MISC ------------------------------------------------------               
        .DMONITOR_CFG                   (24'h000B01),                           // 
        .RX_DEBUG_CFG                   (14'h0000),                             // Optimized for IES
      //.TST_RSV                        (32'd0),                                //
      //.UCODEER_CLR                    ( 1'd0)                                 // 
      
        //---------- GTP -------------------------------------------------------
      //.ACJTAG_DEBUG_MODE              (1'd0),                                 //
      //.ACJTAG_MODE                    (1'd0),                                 //
      //.ACJTAG_RESET                   (1'd0),                                 //
      //.ADAPT_CFG0                     (20'd0),                                //
        .CFOK_CFG                       (43'h490_0004_0E80),                    // Changed from 42 to 43-bits, Optimized for IES
        .CFOK_CFG2                      ( 7'b010_0000),                         // Changed from 6 to 7-bits, Optimized for IES
        .CFOK_CFG3                      ( 7'b010_0000),                         // Changed from 6 to 7-bits, Optimized for IES
        .CFOK_CFG4                      ( 1'd0),                                // GTP new, Optimized for IES
        .CFOK_CFG5                      ( 2'd0),                                // GTP new, Optimized for IES
        .CFOK_CFG6                      ( 4'd0)                                 // GTP new, Optimized for IES
      
     )                                                                        
     model_ap2_tst_gtpe2_channel_i                                                                     
     (                                                                           
                                                                                 
        //---------- Clock -----------------------------------------------------                
        .PLL0CLK                        (GT_QPLLCLK),                           //
        .PLL1CLK                        (1'd0),                                 //
        .PLL0REFCLK                     (GT_QPLLREFCLK),                        //
        .PLL1REFCLK                     (1'd0),                                 //
        .TXUSRCLK                       (GT_TXUSRCLK),                          //
        .RXUSRCLK                       (GT_RXUSRCLK),                          //
        .TXUSRCLK2                      (GT_TXUSRCLK2),                         //
        .RXUSRCLK2                      (GT_RXUSRCLK2),                         //
        .TXSYSCLKSEL                    (GT_TXSYSCLKSEL),                       // 
        .RXSYSCLKSEL                    (GT_RXSYSCLKSEL),                       // 
        .TXOUTCLKSEL                    (txoutclksel),                          //
        .RXOUTCLKSEL                    (rxoutclksel),                          //
        .CLKRSVD0                       (1'd0),                                 // 
        .CLKRSVD1                       (1'd0),                                 // 
                                                                                
        .TXOUTCLK                       (GT_TXOUTCLK),                          //
        .RXOUTCLK                       (GT_RXOUTCLK),                          //
        .TXOUTCLKFABRIC                 (),                                     //
        .RXOUTCLKFABRIC                 (),                                     //
        .TXOUTCLKPCS                    (),                                     //
        .RXOUTCLKPCS                    (),                                     //
        .RXCDRLOCK                      (GT_RXCDRLOCK),                         //
                                                                                
        //---------- Reset -----------------------------------------------------                
        .TXUSERRDY                      (GT_TXUSERRDY),                         //
        .RXUSERRDY                      (GT_RXUSERRDY),                         //
        .CFGRESET                       (1'd0),                                 //
        .GTRESETSEL                     (1'd0),                                 //
        .RESETOVRD                      (GT_RESETOVRD),                         //
        .GTTXRESET                      (GT_GTTXRESET),                         //
        .GTRXRESET                      (GT_GTRXRESET),                         //
                                                                               
        .TXRESETDONE                    (GT_TXRESETDONE),                       //
        .RXRESETDONE                    (GT_RXRESETDONE),                       //
                                                                                
        //---------- TX Data ---------------------------------------------------                
        .TXDATA                         (GT_TXDATA),                            //
        .TXCHARISK                      (GT_TXDATAK),                           //
                                                                                
        .GTPTXP                         (GT_TXP),                               // GTP
        .GTPTXN                         (GT_TXN),                               // GTP 
                                                                                
        //---------- RX Data ---------------------------------------------------                
        .GTPRXP                         (GT_RXP),                               // GTP 
        .GTPRXN                         (GT_RXN),                               // GTP
                                                                              
        .RXDATA                         (rxdata[31:0]),                         //
        .RXCHARISK                      (rxdatak[3:0]),                         //
                                                                                
        //---------- Command ---------------------------------------------------                
        .TXDETECTRX                     (GT_TXDETECTRX),                        //
        .TXPDELECIDLEMODE               ( 1'd0),                                //
        .RXELECIDLEMODE                 ( 2'd0),                                //
        .TXELECIDLE                     (GT_TXELECIDLE),                        //
        .TXCHARDISPMODE                 ({3'd0, GT_TXCOMPLIANCE}),              // Changed from 8 to 4-bits
        .TXCHARDISPVAL                  ( 4'd0),                                // Changed from 8 to 4-bits
        .TXPOLARITY                     ( 1'b0),                                // 
        .RXPOLARITY                     (GT_RXPOLARITY),                        //
        .TXPD                           (GT_TXPOWERDOWN),                       //
        .RXPD                           (GT_RXPOWERDOWN),                       //
        .TXRATE                         (GT_TXRATE),                            //
        .RXRATE                         (GT_RXRATE),                            //
        .TXRATEMODE                     (1'b0),                                 //
        .RXRATEMODE                     (1'b0),                                 //
                                                                                
        //---------- Electrical Command ----------------------------------------                
        .TXMARGIN                       (GT_TXMARGIN),                          //
        .TXSWING                        (GT_TXSWING),                           //
        .TXDEEMPH                       (GT_TXDEEMPH),                          //
        .TXINHIBIT                      (1'd0),                                 // 
        .TXBUFDIFFCTRL                  (3'b100),                               // 
        .TXDIFFCTRL                     (4'b1100),                              // Select 850mV 
        .TXPRECURSOR                    (GT_TXPRECURSOR),                       // 
        .TXPRECURSORINV                 (1'd0),                                 // 
        .TXMAINCURSOR                   (GT_TXMAINCURSOR),                      // 
        .TXPOSTCURSOR                   (GT_TXPOSTCURSOR),                      // 
        .TXPOSTCURSORINV                (1'd0),                                 // 
                                                                                
        //---------- Status ----------------------------------------------------                
        .RXVALID                        (GT_RXVALID),                           //
        .PHYSTATUS                      (GT_PHYSTATUS),                         //
        .RXELECIDLE                     (GT_RXELECIDLE),                        // 
        .RXSTATUS                       (GT_RXSTATUS),                          //
        .TXRATEDONE                     (GT_TXRATEDONE),                        //
        .RXRATEDONE                     (GT_RXRATEDONE),                        //
                                                                                
        //---------- DRP -------------------------------------------------------                
        .DRPCLK                         (GT_DRPCLK),                            //
        .DRPADDR                        (GT_DRPADDR),                           //
        .DRPEN                          (GT_DRPEN),                             //
        .DRPDI                          (GT_DRPDI),                             //
        .DRPWE                          (GT_DRPWE),                             //
                                                                                
        .DRPDO                          (GT_DRPDO),                             //
        .DRPRDY                         (GT_DRPRDY),                            //
                                                                                
        //---------- PMA -------------------------------------------------------                
        .TXPMARESET                     (GT_TXPMARESET),                        //
        .RXPMARESET                     (GT_RXPMARESET),                        //
        .RXLPMRESET                     ( 1'd0),		                            // GTP new  
        .RXLPMOSINTNTRLEN               ( 1'd0),                                // GTP new   
        .RXLPMHFHOLD                    ( 1'd0),                                // 
        .RXLPMHFOVRDEN                  ( 1'd0),                                // 
        .RXLPMLFHOLD                    ( 1'd0),                                // 
        .RXLPMLFOVRDEN                  ( 1'd0),                                // 
        .PMARSVDIN0                     ( 1'd0),                                // GTP new 
        .PMARSVDIN1                     ( 1'd0),                                // GTP new 
        .PMARSVDIN2                     ( 1'd0),                                // GTP new  
        .PMARSVDIN3                     ( 1'd0),                                // GTP new 
        .PMARSVDIN4                     ( 1'd0),                                // GTP new 
        .GTRSVD                         (16'd0),                                // 
              
        .PMARSVDOUT0                    (),                                     // GTP new
        .PMARSVDOUT1                    (),                                     // GTP new                                                                       
        .DMONITOROUT                    (dmonitorout),                          // GTP 15-bits 
                                                                              
        //---------- PCS -------------------------------------------------------                
        .TXPCSRESET                     (GT_TXPCSRESET),                        //
        .RXPCSRESET                     (GT_RXPCSRESET),                        //
        .PCSRSVDIN                      (16'd0),                                // [0]: 1 = TXRATE async, [1]: 1 = RXRATE async    
        
        .PCSRSVDOUT                     (),                                     // 
        
        //---------- CDR -------------------------------------------------------                
        .RXCDRRESET                     (GT_RXCDRRESET),                        //
        .RXCDRRESETRSV                  (1'd0),                                 // 
        .RXCDRFREQRESET                 (GT_RXCDRFREQRESET),                    // 
        .RXCDRHOLD                      (1'b0),                                 //
        .RXCDROVRDEN                    (1'd0),                                 // 
         
        //---------- PI --------------------------------------------------------
        .TXPIPPMEN                      (1'd0),                                 //
        .TXPIPPMOVRDEN                  (1'd0),                                 //
        .TXPIPPMPD                      (1'd0),                                 //
        .TXPIPPMSEL                     (1'd0),                                 //
        .TXPIPPMSTEPSIZE                (5'd0),                                 // 
        .TXPISOPD                       (1'd0),                                 // GTP new 
         
        //---------- DFE -------------------------------------------------------                
        .RXDFEXYDEN                     (1'd0),                                 //  
        
        //---------- OS --------------------------------------------------------         
        .RXOSHOLD                       (1'd0),                                 // Optimized for IES
        .RXOSOVRDEN                     (1'd0),                                 // Optimized for IES                          
        .RXOSINTEN                      (1'd1),                                 // Optimized for IES           
        .RXOSINTHOLD                    (1'd0),                                 // Optimized for IES                                                                                                      
        .RXOSINTNTRLEN                  (1'd0),                                 // Optimized for IES           
        .RXOSINTOVRDEN                  (1'd0),                                 // Optimized for IES            
        .RXOSINTPD                      (1'd0),                                 // GTP new, Optimized for IES             
        .RXOSINTSTROBE                  (1'd0),                                 // Optimized for IES           
        .RXOSINTTESTOVRDEN              (1'd0),                                 // Optimized for IES           
        .RXOSINTCFG                     (4'b0010),                              // Optimized for IES                     
        .RXOSINTID0                     (4'd0),                                 // Optimized for IES
                                  
        .RXOSINTDONE                    (),                                     //
        .RXOSINTSTARTED                 (),                                     //
        .RXOSINTSTROBEDONE              (),                                     //
        .RXOSINTSTROBESTARTED           (),                                     //
                                                                                
        //---------- Eye Scan --------------------------------------------------                
        .EYESCANRESET                   (GT_EYESCANRESET),                      // 
        .EYESCANMODE                    (1'd0),                                 // 
        .EYESCANTRIGGER                 (1'b0),                                 // 
                                                                                
        .EYESCANDATAERROR               (GT_EYESCANDATAERROR),                  //
                                                                                
        //---------- TX Buffer -------------------------------------------------                
        .TXBUFSTATUS                    (),                                     //
                                                                                
        //---------- RX Buffer -------------------------------------------------                
        .RXBUFRESET                     (GT_RXBUFRESET),                        // 
        
        .RXBUFSTATUS                    (GT_RXBUFSTATUS),                       //
                                                                                
        //---------- TX Sync ---------------------------------------------------                
        .TXPHDLYRESET                   (GT_TXPHDLYRESET),                      //
        .TXPHDLYTSTCLK                  (1'd0),                                 //
        .TXPHALIGN                      (GT_TXPHALIGN),                         // 
        .TXPHALIGNEN                    (GT_TXPHALIGNEN),                       //  
        .TXPHDLYPD                      (1'd0),                                 // 
        .TXPHINIT                       (GT_TXPHINIT),                          //  
        .TXPHOVRDEN                     (1'd0),                                 //
        .TXDLYBYPASS                    (GT_TXDLYBYPASS),                       //  
        .TXDLYSRESET                    (GT_TXDLYSRESET),                       // 
        .TXDLYEN                        (GT_TXDLYEN),                           //  
        .TXDLYOVRDEN                    (1'd0),                                 //
        .TXDLYHOLD                      (1'd0),                                 // 
        .TXDLYUPDOWN                    (1'd0),                                 //
                                                                                
        .TXPHALIGNDONE                  (GT_TXPHALIGNDONE),                     // 
        .TXPHINITDONE                   (GT_TXPHINITDONE),                      // 
        .TXDLYSRESETDONE                (GT_TXDLYSRESETDONE),                   //
        
        .TXSYNCMODE                     (GT_TXSYNCMODE),                        //
        .TXSYNCIN                       (GT_TXSYNCIN),                          //
        .TXSYNCALLIN                    (GT_TXSYNCALLIN),                       //
        
        .TXSYNCDONE                     (GT_TXSYNCDONE),                        //
        .TXSYNCOUT                      (GT_TXSYNCOUT),                         //
        
        //---------- RX Sync ---------------------------------------------------                  
        .RXPHDLYRESET                   (1'd0),                                 //
        .RXPHALIGN                      (GT_RXPHALIGN),                         //
        .RXPHALIGNEN                    (GT_RXPHALIGNEN),                       //
        .RXPHDLYPD                      (1'd0),                                 // 
        .RXPHOVRDEN                     (1'd0),                                 // 
        .RXDLYBYPASS                    (GT_RXDLYBYPASS),                       //  
        .RXDLYSRESET                    (GT_RXDLYSRESET),                       // 
        .RXDLYEN                        (GT_RXDLYEN),                           // 
        .RXDLYOVRDEN                    (1'd0),                                 //
        .RXDDIEN                        (GT_RXDDIEN),                           //
                                                                                
        .RXPHALIGNDONE                  (GT_RXPHALIGNDONE),                     //  
        .RXPHMONITOR                    (),                                     //
        .RXPHSLIPMONITOR                (),                                     // 
        .RXDLYSRESETDONE                (GT_RXDLYSRESETDONE),                   // 

        .RXSYNCMODE                     (GT_RXSYNCMODE),                        //
        .RXSYNCIN                       (GT_RXSYNCIN),                          //
        .RXSYNCALLIN                    (GT_RXSYNCALLIN),                       //
        
        .RXSYNCDONE                     (GT_RXSYNCDONE),                        //
        .RXSYNCOUT                      (GT_RXSYNCOUT),                         //
                
        //---------- Comma Alignment -------------------------------------------                 
        .RXCOMMADETEN                   (1'd1),                                 //
        .RXMCOMMAALIGNEN                (1'd1),                                 // No Gen3 support in GTP
        .RXPCOMMAALIGNEN                (1'd1),                                 // No Gen3 support in GTP
        .RXSLIDE                        (GT_RXSLIDE),                           //
        .RXCOMMADET                     (GT_RXCOMMADET),                        //
        .RXCHARISCOMMA                  (rxchariscomma[3:0]),                   // 
        .RXBYTEISALIGNED                (GT_RXBYTEISALIGNED),                   //
        .RXBYTEREALIGN                  (GT_RXBYTEREALIGN),                     //
                                                                                
        //---------- Channel Bonding -------------------------------------------                
        .RXCHBONDEN                     (GT_RXCHBONDEN),                        //
        .RXCHBONDI                      (GT_RXCHBONDI[3:0]),                    //
        .RXCHBONDLEVEL                  (GT_RXCHBONDLEVEL),                     //
        .RXCHBONDMASTER                 (GT_RXCHBONDMASTER),                    //
        .RXCHBONDSLAVE                  (GT_RXCHBONDSLAVE),                     //
                                                                                
        .RXCHANBONDSEQ                  (),                                     // 
        .RXCHANISALIGNED                (GT_RXCHANISALIGNED),                   //
        .RXCHANREALIGN                  (),                                     //
        .RXCHBONDO                      (GT_RXCHBONDO[3:0]),                    //
                                                                                
        //---------- Clock Correction  -----------------------------------------                
        .RXCLKCORCNT                    (),                                     //
                                                                                
        //---------- 8b10b -----------------------------------------------------                
        .TX8B10BBYPASS                  (4'd0),                                 //
        .TX8B10BEN                      (1'b1),                                 // No Gen3 support in GTP
        .RX8B10BEN                      (1'b1),                                 // No Gen3 support in GTP
                                                                                
        .RXDISPERR                      (GT_RXDISPERR[3:0]),                         //
        .RXNOTINTABLE                   (GT_RXNOTINTABLE[3:0]),                      //
                                                                                
        //---------- 64b/66b & 64b/67b -----------------------------------------                  
        .TXHEADER                       (3'd0),                                 //
        .TXSEQUENCE                     (7'd0),                                 //
        .TXSTARTSEQ                     (1'd0),                                 //                                                              
        .RXGEARBOXSLIP                  (1'd0),                                 //
                                                                                
        .TXGEARBOXREADY                 (),                                     // 
        .RXDATAVALID                    (),                                     //
        .RXHEADER                       (),                                     //
        .RXHEADERVALID                  (),                                     //
        .RXSTARTOFSEQ                   (),                                     //
                                                                                
        //---------- PRBS/Loopback ---------------------------------------------                
        .TXPRBSSEL                      (GT_TXPRBSSEL),                         //
        .RXPRBSSEL                      (GT_RXPRBSSEL),                         //
        .TXPRBSFORCEERR                 (GT_TXPRBSFORCEERR),                    //
        .RXPRBSCNTRESET                 (GT_RXPRBSCNTRESET),                    // 
        .LOOPBACK                       (GT_LOOPBACK),                          // 
                                                                                
        .RXPRBSERR                      (GT_RXPRBSERR),                         //
                                                                                
        //---------- OOB -------------------------------------------------------      
        .SIGVALIDCLK                    (GT_OOBCLK),                            // Optimized for debug           
        .TXCOMINIT                      (1'd0),                                 //
        .TXCOMSAS                       (1'd0),                                 //
        .TXCOMWAKE                      (1'd0),                                 //
        .RXOOBRESET                     (1'd0),                                 // 
                                                                                
        .TXCOMFINISH                    (),                                     //
        .RXCOMINITDET                   (),                                     //
        .RXCOMSASDET                    (),                                     //
        .RXCOMWAKEDET                   (),                                     //
                                                                                
        //---------- MISC ------------------------------------------------------                
        .SETERRSTATUS                   ( 1'd0),                                // 
        .TXDIFFPD                       ( 1'd0),                                // 
        .TSTIN                          (20'hFFFFF),                            //  
                 
        //---------- GTP -------------------------------------------------------                                                                        
        .RXADAPTSELTEST                 (14'd0),                                //
        .DMONFIFORESET                  ( 1'd0),                                //
        .DMONITORCLK                    (dmonitorclk),                          //  
        .RXOSCALRESET                   ( 1'd0),                                //                     
                             
        .RXPMARESETDONE                 (GT_RXPMARESETDONE),                    // GTP
        .TXPMARESETDONE                 ()                                      //
        
     );         
     
     assign GT_CPLLLOCK = 1'b0;

    end

else if (PCIE_GT_DEVICE == "GTH") 

    begin : gth_channel
    
    //---------- GTH Channel Module --------------------------------------------
    GTHE2_CHANNEL #
    (
               
        //---------- Simulation Attributes -------------------------------------               
        .SIM_CPLLREFCLK_SEL             (3'b001),                               //
        .SIM_RESET_SPEEDUP              (PCIE_SIM_SPEEDUP),                     //
        .SIM_RECEIVER_DETECT_PASS       ("TRUE"),                               //    
        .SIM_TX_EIDLE_DRIVE_LEVEL       (PCIE_SIM_TX_EIDLE_DRIVE_LEVEL),        // 
        .SIM_VERSION                    ("2.0"),                                //
                                                                               
        //---------- Clock Attributes ------------------------------------------                                      
        .CPLL_REFCLK_DIV                (CPLL_REFCLK_DIV),                      //
        .CPLL_FBDIV_45                  (CPLL_FBDIV_45),                        //
        .CPLL_FBDIV                     (CPLL_FBDIV),                           //
        .TXOUT_DIV                      (OUT_DIV),                              //
        .RXOUT_DIV                      (OUT_DIV),                              // 
        .TX_CLK25_DIV                   (CLK25_DIV),                            //
        .RX_CLK25_DIV                   (CLK25_DIV),                            //
        .TX_CLKMUX_PD                   ( 1'b1),                                // GTH
        .RX_CLKMUX_PD                   ( 1'b1),                                // GTH
        .TX_XCLK_SEL                    (TX_XCLK_SEL),                          // TXOUT = use TX buffer, TXUSR = bypass TX buffer
        .RX_XCLK_SEL                    ("RXREC"),                              // RXREC = use RX buffer, RXUSR = bypass RX buffer
        .OUTREFCLK_SEL_INV              ( 2'b11),                               //
        .CPLL_CFG                       (29'h00A407CC),                         // Changed from 24 to 29-bits, Optimized for PCIe PLL BW 
        .CPLL_INIT_CFG                  (24'h00001E),                           // Optimized for IES
        .CPLL_LOCK_CFG                  (16'h01E8),                             // Optimized for IES
      //.USE_PCS_CLK_PHASE_SEL          ( 1'd0)                                 // GTH new
                                                                               
        //---------- Reset Attributes ------------------------------------------                
        .TXPCSRESET_TIME                (5'b00001),                             //
        .RXPCSRESET_TIME                (5'b00001),                             //
        .TXPMARESET_TIME                (5'b00011),                             //
        .RXPMARESET_TIME                (5'b00011),                             // Optimized for sim and for DRP
      //.RXISCANRESET_TIME              (5'b00001),                             //
      //.RESET_POWERSAVE_DISABLE        ( 1'd0),                                // GTH new
                                                                               
        //---------- TX Data Attributes ----------------------------------------                
        .TX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        .TX_INT_DATAWIDTH               ( 0),                                   // 2-byte internal datawidth for Gen1/Gen2
                                                                               
        //---------- RX Data Attributes ----------------------------------------                
        .RX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        .RX_INT_DATAWIDTH               ( 0),                                   // 2-byte internal datawidth for Gen1/Gen2
                                                                               
        //---------- Command Attributes ----------------------------------------                
        .TX_RXDETECT_CFG                (TX_RXDETECT_CFG),                      //
        .TX_RXDETECT_PRECHARGE_TIME     (17'h00001),                            // GTH new, Optimized for sim
        .TX_RXDETECT_REF                ( 3'b011),                              // 
        .RX_CM_SEL                      ( 2'b11),                                // 0 = AVTT, 1 = GND, 2 = Float, 3 = Programmable, optimized for silicon
        .RX_CM_TRIM                     ( 4'b1010),                             // Select 800mV, Changed from 3 to 4-bits, optimized for silicon
        .TX_EIDLE_ASSERT_DELAY          (PCIE_TX_EIDLE_ASSERT_DELAY),           // Optimized for sim (3'd4)
        .TX_EIDLE_DEASSERT_DELAY        ( 3'b100),                              // Optimized for sim
      //.PD_TRANS_TIME_FROM_P2          (12'h03C),                              //
        .PD_TRANS_TIME_NONE_P2          ( 8'h09),                               // Optimized for sim
      //.PD_TRANS_TIME_TO_P2            ( 8'h64),                               //
      //.TRANS_TIME_RATE                ( 8'h0E),                               //
                                                                               
        //---------- Electrical Command Attributes -----------------------------                
        .TX_DRIVE_MODE                  ("PIPE"),                               // Gen1/Gen2 = PIPE, Gen3 = PIPEGEN3
        .TX_DEEMPH0                     ( 6'b010100),                           //  6.0 dB, optimized for compliance, changed from 5 to 6-bits
        .TX_DEEMPH1                     ( 6'b001011),                           //  3.5 dB, optimized for compliance, changed from 5 to 6-bits
        .TX_MARGIN_FULL_0               ( 7'b1001111),                          // 1000 mV
        .TX_MARGIN_FULL_1               ( 7'b1001110),                          //  950 mV
        .TX_MARGIN_FULL_2               ( 7'b1001101),                          //  900 mV
        .TX_MARGIN_FULL_3               ( 7'b1001100),                          //  850 mV
        .TX_MARGIN_FULL_4               ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_0                ( 7'b1000101),                          //  500 mV
        .TX_MARGIN_LOW_1                ( 7'b1000110),                          //  450 mV
        .TX_MARGIN_LOW_2                ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_3                ( 7'b1000010),                          //  350 mV
        .TX_MARGIN_LOW_4                ( 7'b1000000),                          //  250 mV
        .TX_MAINCURSOR_SEL              ( 1'b0),                                //
        .TX_QPI_STATUS_EN               ( 1'b0),                                //
                                                                               
        //---------- Status Attributes -----------------------------------------                
        .RX_SIG_VALID_DLY               (4),                                    // Optimized for sim
                                                                               
        //---------- DRP Attributes --------------------------------------------                
                     
        //---------- PCS Attributes --------------------------------------------                
        .PCS_PCIE_EN                    ("TRUE"),                               // PCIe 
        .PCS_RSVD_ATTR                  (48'h0000_0000_0140),                   // [8] : 1 = OOB power-up, [6] : 1 = DMON enable, Optimized for IES       
                                                                               
        //---------- PMA Attributes --------------------------------------------                
        .PMA_RSV                        (32'h00000080),                         // Optimized for IES 
        .PMA_RSV2                       (32'h1C00000A),                         // Changed from 16 to 32-bits, Optimized for IES
      //.PMA_RSV3                       ( 2'h0),                                // 
        .PMA_RSV4                       (15'h0008),                             // GTH new, Optimized for IES
      //.PMA_RSV5                       ( 4'h00),                               // GTH new
        .RX_BIAS_CFG                    (24'h0C0010),                           // Changed from 12 to 24-bits, Optimized for IES
        .TERM_RCAL_CFG                  (15'b100001000010000),                  // Changed from  5 to 15-bits, Optimized for IES
        .TERM_RCAL_OVRD                 ( 3'b000),                              // Changed from  1 to  3-bits, Optimized for IES
                  
        //---------- TX PI -----------------------------------------------------             
      //.TXPI_CFG0                      ( 2'd0),                                // GTH new
      //.TXPI_CFG1                      ( 2'd0),                                // GTH new
      //.TXPI_CFG2                      ( 2'd0),                                // GTH new
      //.TXPI_CFG3                      ( 1'd0),                                // GTH new
      //.TXPI_CFG4                      ( 1'd0),                                // GTH new
      //.TXPI_CFG5                      ( 3'b100),                              // GTH new 
      //.TXPI_GREY_SEL                  ( 1'd0),                                // GTH new
      //.TXPI_INVSTROBE_SEL             ( 1'd0),                                // GTH new
      //.TXPI_PPMCLK_SEL                ("TXUSRCLK2"),                          // GTH new
      //.TXPI_PPM_CFG                   ( 8'd0),                                // GTH new
      //.TXPI_SYNFREQ_PPM               ( 3'd0),                                // GTH new
              
        //---------- RX PI -----------------------------------------------------  
        .RXPI_CFG0                      (2'b00),                                // GTH new
        .RXPI_CFG1                      (2'b11),                                // GTH new
        .RXPI_CFG2                      (2'b11),                                // GTH new
        .RXPI_CFG3                      (2'b11),                                // GTH new
        .RXPI_CFG4                      (1'b0),                                 // GTH new
        .RXPI_CFG5                      (1'b0),                                 // GTH new
        .RXPI_CFG6                      (3'b100),                               // GTH new

        //---------- CDR Attributes --------------------------------------------
        .RXCDR_CFG                      (RXCDR_CFG_GTH),                        //
      //.RXCDR_CFG                      (83'h0_0011_07FE_4060_0104_1010),       // A. Changed from 72 to 83-bits, optimized for IES div1 (Gen2), +/-000ppm, default, converted from GTX GES VnC,(2 Gen1)
      //.RXCDR_CFG                      (83'h0_0011_07FE_4060_2104_1010),       // B. Changed from 72 to 83-bits, optimized for IES div1 (Gen2), +/-300ppm, default, converted from GTX GES VnC,(2 Gen1)
      //.RXCDR_CFG                      (83'h0_0011_07FE_2060_0104_1010),       // C. Changed from 72 to 83-bits, optimized for IES div1 (Gen2), +/-000ppm, converted from GTX GES recommended, (3 Gen1)
      //.RXCDR_CFG                      (83'h0_0011_07FE_2060_2104_1010),       // D. Changed from 72 to 83-bits, optimized for IES div1 (Gen2), +/-300ppm, converted from GTX GES recommended, (3 Gen1)
      //.RXCDR_CFG                      (83'h0_0001_07FE_1060_0110_1010),       // E. Changed from 72 to 83-bits, optimized for IES div2 (Gen1), +/-000ppm, default, (3 Gen2)
      //.RXCDR_CFG                      (83'h0_0001_07FE_1060_2110_1010),       // F. Changed from 72 to 83-bits, optimized for IES div2 (Gen1), +/-300ppm, default, (3 Gen2)
      //.RXCDR_CFG                      (83'h0_0011_07FE_1060_0110_1010),       // G. Changed from 72 to 83-bits, optimized for IES div2 (Gen1), +/-000ppm, converted from GTX GES recommended, (3 Gen2)
      //.RXCDR_CFG                      (83'h0_0011_07FE_1060_2110_1010),       // H. Changed from 72 to 83-bits, optimized for IES div2 (Gen1), +/-300ppm, converted from GTX GES recommended, (2 Gen1)
        .RXCDR_LOCK_CFG                 ( 6'b010101),                           // [5:3] Window Refresh, [2:1] Window Size, [0] Enable Detection (sensitive lock = 6'b111001)
        .RXCDR_HOLD_DURING_EIDLE        ( 1'd1),                                // Hold  RX CDR           on electrical idle for Gen1/Gen2
        .RXCDR_FR_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR frequency on electrical idle for Gen3
        .RXCDR_PH_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR phase     on electrical idle for Gen3
      //.RXCDRFREQRESET_TIME            ( 5'b00001),                            // optimized for IES
      //.RXCDRPHRESET_TIME              ( 5'b00001),                            // optimized for IES
                         
        //---------- LPM Attributes --------------------------------------------               
        .RXLPM_HF_CFG                   (14'h0200),                             // Optimized for IES   
        .RXLPM_LF_CFG                   (18'h09000),                            // Changed from 14 to 18-bits, Optimized for IES       
                                                                                
        //---------- DFE Attributes --------------------------------------------                
        .RXDFELPMRESET_TIME	            ( 7'h0F),                               // Optimized for IES     
        .RX_DFE_AGC_CFG0                ( 2'h0),                                // GTH new, optimized for IES    
        .RX_DFE_AGC_CFG1                ( 3'h4),                                // GTH new, optimized for IES, DFE
        .RX_DFE_AGC_CFG2                ( 4'h0),                                // GTH new, optimized for IES 
        .RX_DFE_AGC_OVRDEN              ( 1'h1),                                // GTH new, optimized for IES
        .RX_DFE_GAIN_CFG                (23'h0020C0),                           // Optimized for IES
        .RX_DFE_H2_CFG                  (12'h000),                              // Optimized for IES 
        .RX_DFE_H3_CFG                  (12'h040),                              // Optimized for IES
        .RX_DFE_H4_CFG                  (11'h0E0),                              // Optimized for IES
        .RX_DFE_H5_CFG                  (11'h0E0),                              // Optimized for IES
        .RX_DFE_H6_CFG                  (11'h020),                              // GTH new, optimized for IES
        .RX_DFE_H7_CFG                  (11'h020),                              // GTH new, optimized for IES
        .RX_DFE_KL_CFG                  (33'h000000310),                        // Changed from 13 to 33-bits, optimized for IES
        .RX_DFE_KL_LPM_KH_CFG0          ( 2'h2),                                // GTH new, optimized for IES, DFE
        .RX_DFE_KL_LPM_KH_CFG1          ( 3'h2),                                // GTH new, optimized for IES
        .RX_DFE_KL_LPM_KH_CFG2          ( 4'h2),                                // GTH new, optimized for IES
        .RX_DFE_KL_LPM_KH_OVRDEN        ( 1'h1),                                // GTH new, optimized for IES
        .RX_DFE_KL_LPM_KL_CFG0          ( 2'h2),                                // GTH new, optimized for IES, DFE
        .RX_DFE_KL_LPM_KL_CFG1          ( 3'h2),                                // GTH new, optimized for IES
        .RX_DFE_KL_LPM_KL_CFG2          ( 4'h2),                                // GTH new, optimized for IES
        .RX_DFE_KL_LPM_KL_OVRDEN        ( 1'b1),                                // GTH new, optimized for IES
        .RX_DFE_LPM_CFG                 (16'h0080),                             // Optimized for IES  
        .RX_DFELPM_CFG0                 ( 4'h6),                                // GTH new, optimized for IES
        .RX_DFELPM_CFG1                 ( 4'h0),                                // GTH new, optimized for IES
        .RX_DFELPM_KLKH_AGC_STUP_EN     ( 1'h1),                                // GTH new, optimized for IES
        .RX_DFE_LPM_HOLD_DURING_EIDLE   ( 1'h1),                                // PCIe use mode 
        .RX_DFE_ST_CFG                  (54'h00_C100_000C_003F),                // GTH new, optimized for IES
        .RX_DFE_UT_CFG                  (17'h03800),                            // Optimized for IES
        .RX_DFE_VP_CFG                  (17'h03AA3),                            // Optimized for IES
     
        //---------- OS Attributes ---------------------------------------------
        .RX_OS_CFG                      (13'h0080),                             // Optimized for IES
        .A_RXOSCALRESET                 ( 1'd0),                                // GTH new, optimized for IES
        .RXOSCALRESET_TIME              ( 5'b00011),                            // GTH new, optimized for IES
        .RXOSCALRESET_TIMEOUT           ( 5'b00000),                            // GTH new, disable timeout, optimized for IES
      
        //---------- Eye Scan Attributes ---------------------------------------
      //.ES_CLK_PHASE_SEL               ( 1'd0),                                // GTH new
      //.ES_CONTROL                     ( 6'd0),                                //
      //.ES_ERRDET_EN                   ("FALSE"),                              //
        .ES_EYE_SCAN_EN                 ("FALSE"),                               // Optimized for IES
        .ES_HORZ_OFFSET                 (12'h000),                              // Optimized for IES
      //.ES_PMA_CFG                     (10'd0),                                //
      //.ES_PRESCALE                    ( 5'd0),                                //
      //.ES_QUAL_MASK                   (80'd0),                                //
      //.ES_QUALIFIER                   (80'd0),                                //
      //.ES_SDATA_MASK                  (80'd0),                                //
      //.ES_VERT_OFFSET                 ( 9'd0),                                //
                                                                              
        //---------- TX Buffer Attributes --------------------------------------
        .TXBUF_EN                       (PCIE_TXBUF_EN),                        // 
        .TXBUF_RESET_ON_RATE_CHANGE	    ("TRUE"),                               //
                                                                              
        //---------- RX Buffer Attributes --------------------------------------
        .RXBUF_EN                       ("TRUE"),                               //
      //.RX_BUFFER_CFG                  ( 6'd0),                                //
        .RX_DEFER_RESET_BUF_EN          ("TRUE"),                               // 
        .RXBUF_ADDR_MODE                ("FULL"),                               //
        .RXBUF_EIDLE_HI_CNT	            ( 4'd4),                                // Optimized for sim
        .RXBUF_EIDLE_LO_CNT	            ( 4'd0),                                // Optimized for sim
        .RXBUF_RESET_ON_CB_CHANGE       ("TRUE"),                               //
        .RXBUF_RESET_ON_COMMAALIGN      ("FALSE"),                              //
        .RXBUF_RESET_ON_EIDLE           ("TRUE"),                               // PCIe
        .RXBUF_RESET_ON_RATE_CHANGE	    ("TRUE"),                               //
        .RXBUF_THRESH_OVRD              ("FALSE"),                              //
        .RXBUF_THRESH_OVFLW	            (61),                                   //
        .RXBUF_THRESH_UNDFLW            ( 4),                                   //
      //.RXBUFRESET_TIME                ( 5'b00001),                            //
                                                                              
        //---------- TX Sync Attributes ----------------------------------------
      //.TXPH_CFG                       (16'h0780),                             // 
        .TXPH_MONITOR_SEL               ( 5'd0),                                // 
      //.TXPHDLY_CFG                    (24'h084020),                           // [19] : 1 = full range, 0 = half range
      //.TXDLY_CFG                      (16'h001F),                             // 
      //.TXDLY_LCFG	                    ( 9'h030),                              // 
      //.TXDLY_TAP_CFG                  (16'd0),                                // 
        
        .TXSYNC_OVRD                    (TXSYNC_OVRD),                          // GTH new
        .TXSYNC_MULTILANE               (TXSYNC_MULTILANE),                     // GTH new     
        .TXSYNC_SKIP_DA                 (1'b0),                                 // GTH new   
                                                                              
        //---------- RX Sync Attributes ----------------------------------------
      //.RXPH_CFG                       (24'd0),                                //
        .RXPH_MONITOR_SEL               ( 5'd0),                                //
        .RXPHDLY_CFG                    (24'h004020),                           // [19] : 1 = full range, 0 = half range
      //.RXDLY_CFG                      (16'h001F),                             // 
      //.RXDLY_LCFG	                    ( 9'h030),                              // 
      //.RXDLY_TAP_CFG                  (16'd0),                                //
        .RX_DDI_SEL	                    ( 6'd0),                                //
                
        .RXSYNC_OVRD                    (RXSYNC_OVRD),                          // GTH new        
        .RXSYNC_MULTILANE               (RXSYNC_MULTILANE),                     // GTH new    
        .RXSYNC_SKIP_DA                 (1'b0),                                 // GTH new      
                                                                              
        //---------- Comma Alignment Attributes --------------------------------
        .ALIGN_COMMA_DOUBLE             ("FALSE"),                              //   
        .ALIGN_COMMA_ENABLE             (10'b1111111111),                       // PCIe
        .ALIGN_COMMA_WORD               ( 1),                                   //
        .ALIGN_MCOMMA_DET               ("TRUE"),                               //
        .ALIGN_MCOMMA_VALUE             (10'b1010000011),                       //
        .ALIGN_PCOMMA_DET               ("TRUE"),                               //
        .ALIGN_PCOMMA_VALUE             (10'b0101111100),                       //
        .DEC_MCOMMA_DETECT              ("TRUE"),                               //
        .DEC_PCOMMA_DETECT              ("TRUE"),                               //
        .DEC_VALID_COMMA_ONLY           ("FALSE"),                              // PCIe
        .SHOW_REALIGN_COMMA             ("FALSE"),                              // PCIe
        .RXSLIDE_AUTO_WAIT              ( 7),                                   // 
        .RXSLIDE_MODE                   ("PMA"),                                // PCIe
                                                                              
        //---------- Channel Bonding Attributes --------------------------------
        .CHAN_BOND_KEEP_ALIGN           ("TRUE"),                               // PCIe
        .CHAN_BOND_MAX_SKEW             ( 7),                                   // 
        .CHAN_BOND_SEQ_LEN              ( 4),                                   // PCIe
        .CHAN_BOND_SEQ_1_ENABLE         ( 4'b1111),                             //
        .CHAN_BOND_SEQ_1_1              (10'b0001001010),                       // D10.2 (4A) - TS1 
        .CHAN_BOND_SEQ_1_2              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_3              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .CHAN_BOND_SEQ_2_USE            ("TRUE"),                               // PCIe
        .CHAN_BOND_SEQ_2_ENABLE         ( 4'b1111),                             //
        .CHAN_BOND_SEQ_2_1              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_2              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_3              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .FTS_DESKEW_SEQ_ENABLE          ( 4'b1111),                             // 
        .FTS_LANE_DESKEW_EN	            ("TRUE"),                               // PCIe
        .FTS_LANE_DESKEW_CFG            ( 4'b1111),                             // 
                                                                              
        //---------- Clock Correction Attributes -------------------------------
        .CBCC_DATA_SOURCE_SEL           ("DECODED"),                            //
        .CLK_CORRECT_USE                ("TRUE"),                               //
        .CLK_COR_KEEP_IDLE              ("TRUE"),                               // PCIe
        .CLK_COR_MAX_LAT                (CLK_COR_MAX_LAT),                      // 
        .CLK_COR_MIN_LAT                (CLK_COR_MIN_LAT),                      // 
        .CLK_COR_PRECEDENCE             ("TRUE"),                               //
        .CLK_COR_REPEAT_WAIT            ( 0),                                   // 
        .CLK_COR_SEQ_LEN                ( 1),                                   //
        .CLK_COR_SEQ_1_ENABLE           ( 4'b1111),                             //
        .CLK_COR_SEQ_1_1                (10'b0100011100),                       // K28.0 (1C) - SKP
        .CLK_COR_SEQ_1_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_4                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_ENABLE           ( 4'b0000),                             // Disabled
        .CLK_COR_SEQ_2_USE              ("FALSE"),                              //
        .CLK_COR_SEQ_2_1                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_4                (10'b0000000000),                       // Disabled
                                                                              
        //---------- 8b10b Attributes ------------------------------------------
        .RX_DISPERR_SEQ_MATCH           ("TRUE"),                               //
                                                                              
        //---------- 64b/66b & 64b/67b Attributes ------------------------------
        .GEARBOX_MODE                   (3'd0),                                 //
        .TXGEARBOX_EN                   ("FALSE"),                              //
        .RXGEARBOX_EN                   ("FALSE"),                              //
                                                                              
        //---------- PRBS & Loopback Attributes --------------------------------
        .LOOPBACK_CFG                   ( 1'd1),                                // GTH new, enable latch when bypassing TX buffer, equivalent to GTX PCS_RSVD_ATTR[0]
        .RXPRBS_ERR_LOOPBACK            ( 1'd0),                                //
        .TX_LOOPBACK_DRIVE_HIZ          ("FALSE"),                              //
                                                                              
        //---------- OOB & SATA Attributes -------------------------------------
        .TXOOB_CFG                      ( 1'd1),                                // GTH new, filter stale TX data when exiting TX electrical idle, equivalent to GTX PCS_RSVD_ATTR[7]
      //.RXOOB_CFG                      ( 7'b0000110),                          //
        .RXOOB_CLK_CFG                  (RXOOB_CLK_CFG),                        // GTH new
      //.SAS_MAX_COM                    (64),                                   //
      //.SAS_MIN_COM                    (36),                                   //
      //.SATA_BURST_SEQ_LEN             ( 4'b1111),                             //
      //.SATA_BURST_VAL                 ( 3'b100),                              //
      //.SATA_CPLL_CFG                  ("VCO_3000MHZ"),                        //
      //.SATA_EIDLE_VAL                 ( 3'b100),                              //
      //.SATA_MAX_BURST                 ( 8),                                   //
      //.SATA_MAX_INIT                  (21),                                   //
      //.SATA_MAX_WAKE                  ( 7),                                   //
      //.SATA_MIN_BURST                 ( 4),                                   //
      //.SATA_MIN_INIT                  (12),                                   //
      //.SATA_MIN_WAKE                  ( 4),                                   //  
                                                                              
        //---------- MISC ------------------------------------------------------
        .DMONITOR_CFG                   (24'h000AB1),                           // Optimized for debug; [7:4] : 1011 = AGC
      //.DMONITOR_CFG                   (24'h000AB1),                           // Optimized for debug; [7:4] : 0000 = CDR FSM
        .RX_DEBUG_CFG                   (14'b00000011000000),                   // Changed from 12 to 14-bits, optimized for IES
      //.TST_RSV                        (32'd0),                                //
      //.UCODEER_CLR                    ( 1'd0),                                //
        
        //---------- GTH -------------------------------------------------------
      //.ACJTAG_DEBUG_MODE              ( 1'd0),                                // GTH new
      //.ACJTAG_MODE                    ( 1'd0),                                // GTH new
      //.ACJTAG_RESET                   ( 1'd0),                                // GTH new
        .ADAPT_CFG0                     (20'h00C10),                            // GTH new, optimized for IES
        .CFOK_CFG                       (42'h248_0004_0E80),                    // GTH new, optimized for IES, [8] : 1 = Skip CFOK
        .CFOK_CFG2                      ( 6'b100000),                           // GTH new, optimized for IES
        .CFOK_CFG3                      ( 6'b100000)                            // GTH new, optimized for IES
            
    ) 
    model_ap2_tst_gthe2_channel_i 
    (
           
        //---------- Clock -----------------------------------------------------
        .GTGREFCLK                      (1'd0),                                 //
        .GTREFCLK0                      (GT_GTREFCLK0),                         //
        .GTREFCLK1                      (1'd0),                                 //
        .GTNORTHREFCLK0                 (1'd0),                                 //
        .GTNORTHREFCLK1                 (1'd0),                                 //
        .GTSOUTHREFCLK0                 (1'd0),                                 //
        .GTSOUTHREFCLK1                 (1'd0),                                 //
        .QPLLCLK                        (GT_QPLLCLK),                           //
        .QPLLREFCLK                     (GT_QPLLREFCLK),                        //
        .TXUSRCLK                       (GT_TXUSRCLK),                          //
        .RXUSRCLK                       (GT_RXUSRCLK),                          //
        .TXUSRCLK2                      (GT_TXUSRCLK2),                         //
        .RXUSRCLK2                      (GT_RXUSRCLK2),                         //
        .TXSYSCLKSEL                    (GT_TXSYSCLKSEL),                       // 
        .RXSYSCLKSEL                    (GT_RXSYSCLKSEL),                       // 
        .TXOUTCLKSEL                    (txoutclksel),                          //
        .RXOUTCLKSEL                    (rxoutclksel),                          //
        .CPLLREFCLKSEL                  (3'd1),                                 //
        .CPLLLOCKDETCLK                 (1'd0),                                 //
        .CPLLLOCKEN                     (1'd1),                                 // 
        .CLKRSVD0                       (1'd0),                                 // GTH
        .CLKRSVD1                       (1'd0),                                 // GTH
        
        .TXOUTCLK                       (GT_TXOUTCLK),                          //
        .RXOUTCLK                       (GT_RXOUTCLK),                          //
        .TXOUTCLKFABRIC                 (),                                     //
        .RXOUTCLKFABRIC                 (),                                     //
        .TXOUTCLKPCS                    (),                                     //
        .RXOUTCLKPCS                    (),                                     //
        .CPLLLOCK                       (GT_CPLLLOCK),                          // 
        .CPLLREFCLKLOST                 (),                                     // 
        .CPLLFBCLKLOST                  (),                                     // 
        .RXCDRLOCK                      (GT_RXCDRLOCK),                         //
        .GTREFCLKMONITOR                (),                                     // 
                                                                                
        //---------- Reset -----------------------------------------------------                 
        .CPLLPD                         (cpllpd | GT_CPLLPD),                   // 
        .CPLLRESET                      (cpllrst | GT_CPLLRESET),               //
        .TXUSERRDY                      (GT_TXUSERRDY),                         //
        .RXUSERRDY                      (GT_RXUSERRDY),                         //
        .CFGRESET                       (1'd0),                                 //
        .GTRESETSEL                     (1'd0),                                 // 
        .RESETOVRD                      (GT_RESETOVRD),                         //
        .GTTXRESET                      (GT_GTTXRESET),                         //
        .GTRXRESET                      (GT_GTRXRESET),                         //
                                                                               
        .TXRESETDONE                    (GT_TXRESETDONE),                       //
        .RXRESETDONE                    (GT_RXRESETDONE),                       //
                                                                                
        //---------- TX Data ---------------------------------------------------                 
        .TXDATA                         ({32'd0, GT_TXDATA}),                   //
        .TXCHARISK                      ({ 4'd0, GT_TXDATAK}),                  //
                                                                                
        .GTHTXP                         (GT_TXP),                               // GTH
        .GTHTXN                         (GT_TXN),                               // GTH
                                                                                
        //---------- RX Data ---------------------------------------------------                 
        .GTHRXP                         (GT_RXP),                               // GTH
        .GTHRXN                         (GT_RXN),                               // GTH
                                                                                
        .RXDATA                         (rxdata),                               //
        .RXCHARISK                      (rxdatak),                              //
        
        //---------- Command ---------------------------------------------------
        .TXDETECTRX                     (GT_TXDETECTRX),                        //
        .TXPDELECIDLEMODE               ( 1'd0),                                //
        .RXELECIDLEMODE                 ( 2'd0),                                //
        .TXELECIDLE                     (GT_TXELECIDLE),                        //
        .TXCHARDISPMODE                 ({7'd0, GT_TXCOMPLIANCE}),              //
        .TXCHARDISPVAL                  ( 8'd0),                                //
        .TXPOLARITY                     ( 1'b0),                                // 
        .RXPOLARITY                     (GT_RXPOLARITY),                        //
        .TXPD                           (GT_TXPOWERDOWN),                       //
        .RXPD                           (GT_RXPOWERDOWN),                       //
        .TXRATE                         (GT_TXRATE),                            //
        .RXRATE                         (GT_RXRATE),                            //
        .TXRATEMODE                     (1'd0),                                 // GTH
        .RXRATEMODE                     (1'd0),                                 // GTH
         
        //---------- Electrical Command ----------------------------------------
        .TXMARGIN                       (GT_TXMARGIN),                          //
        .TXSWING                        (GT_TXSWING),                           //
        .TXDEEMPH                       (GT_TXDEEMPH),                          //
        .TXINHIBIT                      (1'd0),                                 // 
        .TXBUFDIFFCTRL                  (3'b100),                               // 
        .TXDIFFCTRL                     (4'b1111),                              // Select 850mV 
        .TXPRECURSOR                    (GT_TXPRECURSOR),                       // 
        .TXPRECURSORINV                 (1'd0),                                 // 
        .TXMAINCURSOR                   (GT_TXMAINCURSOR),                      // 
        .TXPOSTCURSOR                   (GT_TXPOSTCURSOR),                      // 
        .TXPOSTCURSORINV                (1'd0),                                 // 
                                                                              
        //---------- Status ----------------------------------------------------
        .RXVALID                        (GT_RXVALID),                           //
        .PHYSTATUS                      (GT_PHYSTATUS),                         //
        .RXELECIDLE                     (GT_RXELECIDLE),                        // 
        .RXSTATUS                       (GT_RXSTATUS),                          //
        .TXRATEDONE                     (GT_TXRATEDONE),                        //
        .RXRATEDONE                     (GT_RXRATEDONE),                        //
                                                                              
        //---------- DRP -------------------------------------------------------
        .DRPCLK                         (GT_DRPCLK),                            //
        .DRPADDR                        (GT_DRPADDR),                           //
        .DRPEN                          (GT_DRPEN),                             //
        .DRPDI                          (GT_DRPDI),                             //
        .DRPWE                          (GT_DRPWE),                             //
                                                                             
        .DRPDO                          (GT_DRPDO),                             // 
        .DRPRDY                         (GT_DRPRDY),                            // 
                                                                              
        //---------- PMA -------------------------------------------------------
        .TXPMARESET                     (GT_TXPMARESET),                        //
        .RXPMARESET                     (GT_RXPMARESET),                        //
        .RXLPMEN                        (rxlpmen),                              // ***
        .RXLPMHFHOLD                    (GT_RX_CONVERGE),                       // Set to 1 after convergence
        .RXLPMHFOVRDEN                  ( 1'd0),                                // 
        .RXLPMLFHOLD                    (GT_RX_CONVERGE),                       // Set to 1 after convergence
        .RXLPMLFKLOVRDEN                ( 1'd0),                                // 
        .TXQPIBIASEN                    ( 1'd0),                                // 
        .TXQPISTRONGPDOWN               ( 1'd0),                                // 
        .TXQPIWEAKPUP                   ( 1'd0),                                // 
        .RXQPIEN                        ( 1'd0),                                // Optimized for IES
        .PMARSVDIN                      ( 5'd0),                                // 
        .GTRSVD                         (16'd0),                                // 
                                                                              
        .TXQPISENP                      (),                                     // 
        .TXQPISENN                      (),                                     // 
        .RXQPISENP                      (),                                     // 
        .RXQPISENN                      (),                                     // 
        .DMONITOROUT                    (dmonitorout),                          // GTH 15-bits.
                                                                              
        //---------- PCS -------------------------------------------------------                 
        .TXPCSRESET                     (GT_TXPCSRESET),                        //
        .RXPCSRESET                     (GT_RXPCSRESET),                        //
        .PCSRSVDIN                      (16'd0),                                // [0]: 1 = TXRATE async, [1]: 1 = RXRATE async  
        .PCSRSVDIN2                     ( 5'd0),                                // 
                                                                                
        .PCSRSVDOUT                     (),                                     // 
       
        //---------- CDR -------------------------------------------------------                  
        .RXCDRRESET                     (GT_RXCDRRESET),                        //
        .RXCDRRESETRSV                  (1'd0),                                 // 
        .RXCDRFREQRESET                 (GT_RXCDRFREQRESET),                    // 
        .RXCDRHOLD                      (1'b0),                                 //
        .RXCDROVRDEN                    (1'd0),                                 // 
                      
         //---------- PI --------------------------------------------------------
        .TXPIPPMEN                      (1'd0),                                 // GTH new
        .TXPIPPMOVRDEN                  (1'd0),                                 // GTH new
        .TXPIPPMPD                      (1'd0),                                 // GTH new
        .TXPIPPMSEL                     (1'd0),                                 // GTH new
        .TXPIPPMSTEPSIZE                (5'd0),                                 // GTH new            
                                                                
        //---------- DFE -------------------------------------------------------   
        .RXDFELPMRESET                  (GT_RXDFELPMRESET),                     //  
        .RXDFEAGCTRL                    (5'b10000),                             // GTH new, optimized for IES
        .RXDFECM1EN                     (1'd0),                                 // 
        .RXDFEVSEN                      (1'd0),                                 // 
        .RXDFETAP2HOLD                  (1'd0),                                 // 
        .RXDFETAP2OVRDEN                (1'd0),                                 // 
        .RXDFETAP3HOLD                  (1'd0),                                 // 
        .RXDFETAP3OVRDEN                (1'd0),                                 // 
        .RXDFETAP4HOLD                  (1'd0),                                 // 
        .RXDFETAP4OVRDEN                (1'd0),                                 // 
        .RXDFETAP5HOLD                  (1'd0),                                 // 
        .RXDFETAP5OVRDEN                (1'd0),                                 // 
        .RXDFETAP6HOLD                  (1'd0),                                 // GTH new
        .RXDFETAP6OVRDEN                (1'd0),                                 // GTH new
        .RXDFETAP7HOLD                  (1'd0),                                 // GTH new
        .RXDFETAP7OVRDEN                (1'd0),                                 // GTH new
        .RXDFEAGCHOLD                   (GT_RX_CONVERGE),                       // Set to 1 after convergence
        .RXDFEAGCOVRDEN                 (rxlpmen),                              // 
        .RXDFELFHOLD                    (GT_RX_CONVERGE),                       // Set to 1 after convergence 
        .RXDFELFOVRDEN                  (1'd0),                                 // 
        .RXDFEUTHOLD                    (1'd0),                                 // 
        .RXDFEUTOVRDEN                  (1'd0),                                 // 
        .RXDFEVPHOLD                    (1'd0),                                 // 
        .RXDFEVPOVRDEN                  (1'd0),                                 // 
        .RXDFEXYDEN                     (1'd1),                                 // Optimized for IES 
        .RXMONITORSEL                   (2'd0),                                 //
        .RXDFESLIDETAP                  (5'd0),                                 // GTH new
        .RXDFESLIDETAPID                (6'd0),                                 // GTH new
        .RXDFESLIDETAPHOLD              (1'd0),                                 // GTH new
        .RXDFESLIDETAPOVRDEN            (1'd0),                                 // GTH new
        .RXDFESLIDETAPADAPTEN           (1'd0),                                 // GTH new
        .RXDFESLIDETAPINITOVRDEN        (1'd0),                                 // GTH new
        .RXDFESLIDETAPONLYADAPTEN       (1'd0),                                 // GTH new
        .RXDFESLIDETAPSTROBE            (1'd0),                                 // GTH new
    
        .RXMONITOROUT                   (),                                     // 
        .RXDFESLIDETAPSTARTED           (),                                     // GTH new
        .RXDFESLIDETAPSTROBEDONE        (),                                     // GTH new
        .RXDFESLIDETAPSTROBESTARTED     (),                                     // GTH new
        .RXDFESTADAPTDONE               (),                                     // GTH new
        
        //---------- OS --------------------------------------------------------
        .RXOSHOLD                       (1'd0),                                 // optimized for IES
        .RXOSOVRDEN                     (1'd0),                                 // optimized for IES
        .RXOSINTEN                      (1'd1),                                 // GTH new, optimized for IES
        .RXOSINTHOLD                    (1'd0),                                 // GTH new, optimized for IES
        .RXOSINTNTRLEN                  (1'd0),                                 // GTH new, optimized for IES
        .RXOSINTOVRDEN                  (1'd0),                                 // GTH new, optimized for IES
        .RXOSINTSTROBE                  (1'd0),                                 // GTH new, optimized for IES
        .RXOSINTTESTOVRDEN              (1'd0),                                 // GTH new, optimized for IES
        .RXOSINTCFG                     (4'b0110),                              // GTH new, optimized for IES
        .RXOSINTID0                     (4'b0000),                              // GTH new, optimized for IES
        .RXOSCALRESET                   ( 1'd0),                                // GTH, optimized for IES
        
        .RSOSINTDONE                    (),                                     // GTH new
        .RXOSINTSTARTED                 (),                                     // GTH new
        .RXOSINTSTROBEDONE              (),                                     // GTH new
        .RXOSINTSTROBESTARTED           (),                                     // GTH new
        
        //---------- Eye Scan --------------------------------------------------
        .EYESCANRESET                   (GT_EYESCANRESET),                      // 
        .EYESCANMODE                    (1'd0),                                 // 
        .EYESCANTRIGGER                 (1'b0),                                 // 
        
        .EYESCANDATAERROR               (GT_EYESCANDATAERROR),                  //
     
        //---------- TX Buffer -------------------------------------------------
        .TXBUFSTATUS                    (),                                     //
        
        //---------- RX Buffer -------------------------------------------------
        .RXBUFRESET                     (GT_RXBUFRESET),                        //
        
        .RXBUFSTATUS                    (GT_RXBUFSTATUS),                       //
       
        //---------- TX Sync ---------------------------------------------------
        .TXPHDLYRESET                   (GT_TXPHDLYRESET),                      //
        .TXPHDLYTSTCLK                  (1'd0),                                 //
        .TXPHALIGN                      (GT_TXPHALIGN),                         // 
        .TXPHALIGNEN                    (GT_TXPHALIGNEN),                       //  
        .TXPHDLYPD                      (1'd0),                                 // 
        .TXPHINIT                       (GT_TXPHINIT),                          //  
        .TXPHOVRDEN                     (1'd0),                                 //
        .TXDLYBYPASS                    (GT_TXDLYBYPASS),                       //  
        .TXDLYSRESET                    (GT_TXDLYSRESET),                       // 
        .TXDLYEN                        (GT_TXDLYEN),                           //  
        .TXDLYOVRDEN                    (1'd0),                                 //
        .TXDLYHOLD                      (1'd0),                                 // 
        .TXDLYUPDOWN                    (1'd0),                                 //
        
        .TXPHALIGNDONE                  (GT_TXPHALIGNDONE),                     // 
        .TXPHINITDONE                   (GT_TXPHINITDONE),                      // 
        .TXDLYSRESETDONE                (GT_TXDLYSRESETDONE),                   //

        .TXSYNCMODE                     (GT_TXSYNCMODE),                        // GTH
        .TXSYNCIN                       (GT_TXSYNCIN),                          // GTH
        .TXSYNCALLIN                    (GT_TXSYNCALLIN),                       // GTH
        
        .TXSYNCDONE                     (GT_TXSYNCDONE),                        // GTH
        .TXSYNCOUT                      (GT_TXSYNCOUT),                         // GTH
        
        //---------- RX Sync ---------------------------------------------------  
        .RXPHDLYRESET                   (1'd0),                                 //
        .RXPHALIGN                      (GT_RXPHALIGN),                         //
        .RXPHALIGNEN                    (GT_RXPHALIGNEN),                       //
        .RXPHDLYPD                      (1'd0),                                 // 
        .RXPHOVRDEN                     (1'd0),                                 // 
        .RXDLYBYPASS                    (GT_RXDLYBYPASS),                       //  
        .RXDLYSRESET                    (GT_RXDLYSRESET),                       // 
        .RXDLYEN                        (GT_RXDLYEN),                           // 
        .RXDLYOVRDEN                    (1'd0),                                 //
        .RXDDIEN                        (GT_RXDDIEN),                           //
        
        .RXPHALIGNDONE                  (GT_RXPHALIGNDONE),                     //  
        .RXPHMONITOR                    (),                                     //
        .RXPHSLIPMONITOR                (),                                     // 
        .RXDLYSRESETDONE                (GT_RXDLYSRESETDONE),                   // 
         
        .RXSYNCMODE                     (GT_RXSYNCMODE),                        // GTH
        .RXSYNCIN                       (GT_RXSYNCIN),                          // GTH
        .RXSYNCALLIN                    (GT_RXSYNCALLIN),                       // GTH
        
        .RXSYNCDONE                     (GT_RXSYNCDONE),                        // GTH
        .RXSYNCOUT                      (GT_RXSYNCOUT),                         // GTH
         
        //---------- Comma Alignment ------------------------------------------- 
        .RXCOMMADETEN                   ( 1'd1),                                //
        .RXMCOMMAALIGNEN                (!GT_GEN3),                             // 0 = disable comma alignment in Gen3
        .RXPCOMMAALIGNEN                (!GT_GEN3),                             // 0 = disable comma alignment in Gen3
        .RXSLIDE                        ( GT_RXSLIDE),                          //
         
        .RXCOMMADET                     (GT_RXCOMMADET),                        //
        .RXCHARISCOMMA                  (rxchariscomma),                        // 
        .RXBYTEISALIGNED                (GT_RXBYTEISALIGNED),                   //
        .RXBYTEREALIGN                  (GT_RXBYTEREALIGN),                     //
         
        //---------- Channel Bonding -------------------------------------------
        .RXCHBONDEN                     (GT_RXCHBONDEN),                        //
        .RXCHBONDI                      (GT_RXCHBONDI),                         //
        .RXCHBONDLEVEL                  (GT_RXCHBONDLEVEL),                     //
        .RXCHBONDMASTER                 (GT_RXCHBONDMASTER),                    //
        .RXCHBONDSLAVE                  (GT_RXCHBONDSLAVE),                     //
    
        .RXCHANBONDSEQ                  (),                                     //
        .RXCHANISALIGNED                (GT_RXCHANISALIGNED),                   //
        .RXCHANREALIGN                  (),                                     //
        .RXCHBONDO                      (GT_RXCHBONDO),                         //
         
        //---------- Clock Correction  -----------------------------------------
        .RXCLKCORCNT                    (),                                     //
         
        //---------- 8b10b -----------------------------------------------------
        .TX8B10BBYPASS                  (8'd0),                                 //
        .TX8B10BEN                      (!GT_GEN3),                             // 0 = disable TX 8b10b in Gen3
        .RX8B10BEN                      (!GT_GEN3),                             // 0 = disable RX 8b10b in Gen3
        
        .RXDISPERR                      (GT_RXDISPERR),                         //
        .RXNOTINTABLE                   (GT_RXNOTINTABLE),                      //
    
        //---------- 64b/66b & 64b/67b -----------------------------------------
        .TXHEADER                       (3'd0),                                 //
        .TXSEQUENCE                     (7'd0),                                 //
        .TXSTARTSEQ                     (1'd0),                                 //
        .RXGEARBOXSLIP                  (1'd0),                                 //
        
        .TXGEARBOXREADY                 (),                                     // 
        .RXDATAVALID                    (),                                     //
        .RXHEADER                       (),                                     //
        .RXHEADERVALID                  (),                                     //
        .RXSTARTOFSEQ                   (),                                     //
        
        //---------- PRBS & Loopback -------------------------------------------
        .TXPRBSSEL                      (GT_TXPRBSSEL),                         //
        .RXPRBSSEL                      (GT_RXPRBSSEL),                         //
        .TXPRBSFORCEERR                 (GT_TXPRBSFORCEERR),                    //
        .RXPRBSCNTRESET                 (GT_RXPRBSCNTRESET),                    // 
        .LOOPBACK                       (GT_LOOPBACK),                          // 
                                                                                
        .RXPRBSERR                      (GT_RXPRBSERR),                         //
         
        //---------- OOB -------------------------------------------------------
        .SIGVALIDCLK                    (GT_OOBCLK),                            // GTH, optimized for debug
        .TXCOMINIT                      (1'd0),                                 //
        .TXCOMSAS                       (1'd0),                                 //
        .TXCOMWAKE                      (1'd0),                                 //
        .RXOOBRESET                     (1'd0),                                 // 
    
        .TXCOMFINISH                    (),                                     //
        .RXCOMINITDET                   (),                                     //
        .RXCOMSASDET                    (),                                     //
        .RXCOMWAKEDET                   (),                                     //
    
        //---------- MISC ------------------------------------------------------
        .SETERRSTATUS                   ( 1'd0),                                // 
        .TXDIFFPD                       ( 1'd0),                                // 
        .TXPISOPD                       ( 1'd0),                                // 
        .TSTIN                          (20'hFFFFF),                            //  
        
        //---------- GTH -------------------------------------------------------
        .RXADAPTSELTEST                 (14'd0),                                // GTH new
        .DMONFIFORESET                  ( 1'd0),                                // GTH
        .DMONITORCLK                    (dmonitorclk),                          // GTH, optimized for debug
      //.DMONITORCLK                    (GT_DRPCLK),                            // GTH, optimized for debug
        
        .RXPMARESETDONE                 (GT_RXPMARESETDONE),                    // GTH
        .TXPMARESETDONE                 ()                                      // GTH

    );
    
    end
    
else

    begin : gtx_channel

    //---------- GTX Channel Module --------------------------------------------
    GTXE2_CHANNEL #
    (
               
        //---------- Simulation Attributes -------------------------------------
        .SIM_CPLLREFCLK_SEL             (3'b001),                               //
        .SIM_RESET_SPEEDUP              (PCIE_SIM_SPEEDUP),                     //
        .SIM_RECEIVER_DETECT_PASS       ("TRUE"),                               //    
        .SIM_TX_EIDLE_DRIVE_LEVEL       (PCIE_SIM_TX_EIDLE_DRIVE_LEVEL),        // 
        .SIM_VERSION                    (PCIE_USE_MODE),                        //
                                                                                
        //---------- Clock Attributes ------------------------------------------                                      
        .CPLL_REFCLK_DIV                (CPLL_REFCLK_DIV),                      //
        .CPLL_FBDIV_45                  (CPLL_FBDIV_45),                        //
        .CPLL_FBDIV                     (CPLL_FBDIV),                           //
        .TXOUT_DIV                      (OUT_DIV),                              //
        .RXOUT_DIV                      (OUT_DIV),                              // 
        .TX_CLK25_DIV                   (CLK25_DIV),                            //
        .RX_CLK25_DIV                   (CLK25_DIV),                            //
        .TX_CLKMUX_PD                   (CLKMUX_PD),                            // GTX
        .RX_CLKMUX_PD                   (CLKMUX_PD),                            // GTX
        .TX_XCLK_SEL                    (TX_XCLK_SEL),                          // TXOUT = use TX buffer, TXUSR = bypass TX buffer
        .RX_XCLK_SEL                    ("RXREC"),                              // RXREC = use RX buffer, RXUSR = bypass RX buffer
        .OUTREFCLK_SEL_INV              ( 2'b11),                               //
        .CPLL_CFG                       (CPLL_CFG),                             // Optimized for silicon
      //.CPLL_INIT_CFG                  (24'h00001E),                           // 
      //.CPLL_LOCK_CFG                  (16'h01E8),                             //
                                                                                
        //---------- Reset Attributes ------------------------------------------                
        .TXPCSRESET_TIME                (5'b00001),                             //
        .RXPCSRESET_TIME                (5'b00001),                             //
        .TXPMARESET_TIME                (5'b00011),                             //
        .RXPMARESET_TIME                (5'b00011),                             // Optimized for sim and for DRP
      //.RXISCANRESET_TIME              (5'b00001),                             //
                                                                                
        //---------- TX Data Attributes ----------------------------------------                
        .TX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        .TX_INT_DATAWIDTH               ( 0),                                   // 2-byte internal datawidth for Gen1/Gen2
                                                                                
        //---------- RX Data Attributes ----------------------------------------                
        .RX_DATA_WIDTH                  (20),                                   // 2-byte external datawidth for Gen1/Gen2
        .RX_INT_DATAWIDTH               ( 0),                                   // 2-byte internal datawidth for Gen1/Gen2
                                                                                
        //---------- Command Attributes ----------------------------------------                
        .TX_RXDETECT_CFG                (TX_RXDETECT_CFG),                      //
        .TX_RXDETECT_REF                (TX_RXDETECT_REF),                      // 
        .RX_CM_SEL                      ( 2'd3),                                // 0 = AVTT, 1 = GND, 2 = Float, 3 = Programmable
        .RX_CM_TRIM	                    ( 3'b010),                              // Select 800mV
        .TX_EIDLE_ASSERT_DELAY          (PCIE_TX_EIDLE_ASSERT_DELAY),           // Optimized for sim (3'd4)
        .TX_EIDLE_DEASSERT_DELAY        ( 3'b100),                              // Optimized for sim
      //.PD_TRANS_TIME_FROM_P2          (12'h03C),                              //
        .PD_TRANS_TIME_NONE_P2          ( 8'h09),                               //
      //.PD_TRANS_TIME_TO_P2            ( 8'h64),                               //
      //.TRANS_TIME_RATE                ( 8'h0E),                               //
                                                                                
        //---------- Electrical Command Attributes -----------------------------                
        .TX_DRIVE_MODE                  ("PIPE"),                               // Gen1/Gen2 = PIPE, Gen3 = PIPEGEN3
        .TX_DEEMPH0                     ( 5'b10100),                            //  6.0 dB
        .TX_DEEMPH1                     ( 5'b01011),                            //  3.5 dB
        .TX_MARGIN_FULL_0               ( 7'b1001111),                          // 1000 mV
        .TX_MARGIN_FULL_1               ( 7'b1001110),                          //  950 mV
        .TX_MARGIN_FULL_2               ( 7'b1001101),                          //  900 mV
        .TX_MARGIN_FULL_3               ( 7'b1001100),                          //  850 mV
        .TX_MARGIN_FULL_4               ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_0                ( 7'b1000101),                          //  500 mV
        .TX_MARGIN_LOW_1                ( 7'b1000110),                          //  450 mV
        .TX_MARGIN_LOW_2                ( 7'b1000011),                          //  400 mV
        .TX_MARGIN_LOW_3                ( 7'b1000010),                          //  350 mV
        .TX_MARGIN_LOW_4                ( 7'b1000000),                          //  250 mV
        .TX_MAINCURSOR_SEL              ( 1'b0),                                //
        .TX_PREDRIVER_MODE              ( 1'b0),                                // GTX
        .TX_QPI_STATUS_EN               ( 1'b0),                                //
                                                                                
        //---------- Status Attributes -----------------------------------------                
        .RX_SIG_VALID_DLY               (4),                                    // Optimized for sim
                                                                                
        //---------- DRP Attributes --------------------------------------------                
                         
        //---------- PCS Attributes --------------------------------------------                
        .PCS_PCIE_EN                    ("TRUE"),                               // PCIe
        .PCS_RSVD_ATTR                  (PCS_RSVD_ATTR),                        //         
                                                                                
        //---------- PMA Attributes --------------------------------------------                
        .PMA_RSV                        (32'h00018480),                         // Optimized for GES Gen1/Gen2
        .PMA_RSV2                       (16'h2050),                             // Optimized for silicon, [4] RX_CM_TRIM[4], [5] = 1 Enable Eye Scan
      //.PMA_RSV3                       ( 2'd0),                                // 
      //.PMA_RSV4                       (32'd0),                                // GTX 3.0 new
        .RX_BIAS_CFG                    (12'b000000000100),                     // Optimized for GES
      //.TERM_RCAL_CFG                  ( 5'b10000),                            // 
      //.TERM_RCAL_OVRD                 ( 1'd0),                                // 
    
        //---------- CDR Attributes --------------------------------------------
        .RXCDR_CFG                      (RXCDR_CFG_GTX),                        // 
        .RXCDR_LOCK_CFG                 ( 6'b010101),                           // [5:3] Window Refresh, [2:1] Window Size, [0] Enable Detection (sensitive lock = 6'b111001)
        .RXCDR_HOLD_DURING_EIDLE        ( 1'd1),                                // Hold  RX CDR           on electrical idle for Gen1/Gen2
        .RXCDR_FR_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR frequency on electrical idle for Gen3
        .RXCDR_PH_RESET_ON_EIDLE        ( 1'd0),                                // Reset RX CDR phase     on electrical idle for Gen3
      //.RXCDRFREQRESET_TIME            ( 5'b00001),                            // 
      //.RXCDRPHRESET_TIME              ( 5'b00001),                            // 
                                 
        //---------- LPM Attributes --------------------------------------------               
        .RXLPM_HF_CFG                   (14'h00F0),                             // Optimized for silicon
        .RXLPM_LF_CFG                   (14'h00F0),                             // Optimized for silicon
                                                                          
        //---------- DFE Attributes --------------------------------------------                
      //.RXDFELPMRESET_TIME	            ( 7'b0001111),                          // 
        .RX_DFE_GAIN_CFG                (23'h020FEA),                           // Optimized for GES, IES = 23'h001F0A 
        .RX_DFE_H2_CFG                  (12'b000000000000),                     // Optimized for GES
        .RX_DFE_H3_CFG                  (12'b000001000000),                     // Optimized for GES
        .RX_DFE_H4_CFG                  (11'b00011110000),                      // Optimized for GES
        .RX_DFE_H5_CFG                  (11'b00011100000),                      // Optimized for GES
        .RX_DFE_KL_CFG                  (13'b0000011111110),                    // Optimized for GES
        .RX_DFE_KL_CFG2                 (32'h3290D86C),                         // Optimized for GES, GTX new, CTLE 3 3 5, default = 32'h3010D90C
        .RX_DFE_LPM_CFG                 (16'h0954),                             // Optimized for GES
        .RX_DFE_LPM_HOLD_DURING_EIDLE   ( 1'd1),                                // Optimized for PCIe
        .RX_DFE_UT_CFG                  (17'b10001111000000000),                // Optimized for GES, IES = 17'h08F00
        .RX_DFE_VP_CFG                  (17'b00011111100000011),                // Optimized for GES
        .RX_DFE_XYD_CFG                 (13'h0000),                             // Optimized for 4.0
      
        //---------- OS Attributes ---------------------------------------------
        .RX_OS_CFG                      (13'b0000010000000),                    // Optimized for GES
                                                                                
        //---------- Eye Scan Attributes ---------------------------------------                
      //.ES_CONTROL                     ( 6'd0),                                //
      //.ES_ERRDET_EN                   ("FALSE"),                              //
        .ES_EYE_SCAN_EN                 ("FALSE"),                               // 
        .ES_HORZ_OFFSET                 (12'd0),                                //
      //.ES_PMA_CFG                     (10'd0),                                //
      //.ES_PRESCALE                    ( 5'd0),                                //
      //.ES_QUAL_MASK                   (80'd0),                                //
      //.ES_QUALIFIER                   (80'd0),                                //
      //.ES_SDATA_MASK                  (80'd0),                                //
      //.ES_VERT_OFFSET                 ( 9'd0),                                //
                                                                                
        //---------- TX Buffer Attributes --------------------------------------               
        .TXBUF_EN                       (PCIE_TXBUF_EN),                        // 
        .TXBUF_RESET_ON_RATE_CHANGE	    ("TRUE"),                               //
                                                                                
        //---------- RX Buffer Attributes --------------------------------------                
        .RXBUF_EN                       ("TRUE"),                               //
      //.RX_BUFFER_CFG                  ( 6'd0),                                //
        .RX_DEFER_RESET_BUF_EN          ("TRUE"),                               // 
        .RXBUF_ADDR_MODE                ("FULL"),                               //
        .RXBUF_EIDLE_HI_CNT	            ( 4'd4),                                // Optimized for sim
        .RXBUF_EIDLE_LO_CNT	            ( 4'd0),                                // Optimized for sim
        .RXBUF_RESET_ON_CB_CHANGE       ("TRUE"),                               //
        .RXBUF_RESET_ON_COMMAALIGN      ("FALSE"),                              //
        .RXBUF_RESET_ON_EIDLE           ("TRUE"),                               // PCIe
        .RXBUF_RESET_ON_RATE_CHANGE	    ("TRUE"),                               //
        .RXBUF_THRESH_OVRD              ("FALSE"),                              //
        .RXBUF_THRESH_OVFLW	            (61),                                   //
        .RXBUF_THRESH_UNDFLW            ( 4),                                   //
      //.RXBUFRESET_TIME                ( 5'b00001),                            //
                                                                                
        //---------- TX Sync Attributes ----------------------------------------                
      //.TXPH_CFG                       (16'h0780),                             // 
        .TXPH_MONITOR_SEL               ( 5'd0),                                // 
      //.TXPHDLY_CFG                    (24'h084020),                           // 
      //.TXDLY_CFG                      (16'h001F),                             // 
      //.TXDLY_LCFG	                    ( 9'h030),                              // 
      //.TXDLY_TAP_CFG                  (16'd0),                                // 
                                                                                
        //---------- RX Sync Attributes ----------------------------------------            
      //.RXPH_CFG                       (24'd0),                                //
        .RXPH_MONITOR_SEL               ( 5'd0),                                //
        .RXPHDLY_CFG                    (24'h004020),                           // Optimized for sim
      //.RXDLY_CFG                      (16'h001F),                             // 
      //.RXDLY_LCFG	                    ( 9'h030),                              //
      //.RXDLY_TAP_CFG                  (16'd0),                                //
        .RX_DDI_SEL	                    ( 6'd0),                                //
                                                                                
        //---------- Comma Alignment Attributes --------------------------------            
        .ALIGN_COMMA_DOUBLE             ("FALSE"),                              //   
        .ALIGN_COMMA_ENABLE             (10'b1111111111),                       // PCIe
        .ALIGN_COMMA_WORD               ( 1),                                   //
        .ALIGN_MCOMMA_DET               ("TRUE"),                               //
        .ALIGN_MCOMMA_VALUE             (10'b1010000011),                       //
        .ALIGN_PCOMMA_DET               ("TRUE"),                               //
        .ALIGN_PCOMMA_VALUE             (10'b0101111100),                       //
        .DEC_MCOMMA_DETECT              ("TRUE"),                               //
        .DEC_PCOMMA_DETECT              ("TRUE"),                               //
        .DEC_VALID_COMMA_ONLY           ("FALSE"),                              // PCIe
        .SHOW_REALIGN_COMMA             ("FALSE"),                              // PCIe
        .RXSLIDE_AUTO_WAIT              ( 7),                                   // 
        .RXSLIDE_MODE                   ("PMA"),                                // PCIe
                                                                                
        //---------- Channel Bonding Attributes --------------------------------                
        .CHAN_BOND_KEEP_ALIGN           ("TRUE"),                               // PCIe
        .CHAN_BOND_MAX_SKEW             ( 7),                                   // 
        .CHAN_BOND_SEQ_LEN              ( 4),                                   // PCIe
        .CHAN_BOND_SEQ_1_ENABLE         ( 4'b1111),                             //
        .CHAN_BOND_SEQ_1_1              (10'b0001001010),                       // D10.2 (4A) - TS1 
        .CHAN_BOND_SEQ_1_2              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_3              (10'b0001001010),                       // D10.2 (4A) - TS1
        .CHAN_BOND_SEQ_1_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .CHAN_BOND_SEQ_2_USE            ("TRUE"),                               // PCIe
        .CHAN_BOND_SEQ_2_ENABLE         ( 4'b1111),                             //
        .CHAN_BOND_SEQ_2_1              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_2              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_3              (10'b0001000101),                       // D5.2  (45) - TS2
        .CHAN_BOND_SEQ_2_4              (10'b0110111100),                       // K28.5 (BC) - COM
        .FTS_DESKEW_SEQ_ENABLE          ( 4'b1111),                             // 
        .FTS_LANE_DESKEW_EN	            ("TRUE"),                               // PCIe
        .FTS_LANE_DESKEW_CFG            ( 4'b1111),                             // 
                                                                                
        //---------- Clock Correction Attributes -------------------------------            
        .CBCC_DATA_SOURCE_SEL           ("DECODED"),                            //
        .CLK_CORRECT_USE                ("TRUE"),                               //
        .CLK_COR_KEEP_IDLE              ("TRUE"),                               // PCIe
        .CLK_COR_MAX_LAT                (CLK_COR_MAX_LAT),                      // 
        .CLK_COR_MIN_LAT                (CLK_COR_MIN_LAT),                      // 
        .CLK_COR_PRECEDENCE             ("TRUE"),                               //
        .CLK_COR_REPEAT_WAIT            ( 0),                                   // 
        .CLK_COR_SEQ_LEN                ( 1),                                   //
        .CLK_COR_SEQ_1_ENABLE           ( 4'b1111),                             //
        .CLK_COR_SEQ_1_1                (10'b0100011100),                       // K28.0 (1C) - SKP
        .CLK_COR_SEQ_1_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_1_4                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_ENABLE           ( 4'b0000),                             // Disabled
        .CLK_COR_SEQ_2_USE              ("FALSE"),                              //
        .CLK_COR_SEQ_2_1                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_2                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_3                (10'b0000000000),                       // Disabled
        .CLK_COR_SEQ_2_4                (10'b0000000000),                       // Disabled
                                                                                
        //---------- 8b10b Attributes ------------------------------------------                
        .RX_DISPERR_SEQ_MATCH           ("TRUE"),                               //
                                                                                
        //---------- 64b/66b & 64b/67b Attributes ------------------------------                
        .GEARBOX_MODE                   (3'd0),                                 //
        .TXGEARBOX_EN                   ("FALSE"),                              //
        .RXGEARBOX_EN                   ("FALSE"),                              //
                                                                                
        //---------- PRBS & Loopback Attributes --------------------------------                
        .RXPRBS_ERR_LOOPBACK            (1'd0),                                 //
        .TX_LOOPBACK_DRIVE_HIZ          ("FALSE"),                              //
                                                                                
        //---------- OOB & SATA Attributes -------------------------------------                
      //.RXOOB_CFG                      ( 7'b0000110),                          //
      //.SAS_MAX_COM                    (64),                                   //
      //.SAS_MIN_COM                    (36),                                   //
      //.SATA_BURST_SEQ_LEN             ( 4'b1111),                             //
      //.SATA_BURST_VAL                 ( 3'b100),                              //
      //.SATA_CPLL_CFG                  ("VCO_3000MHZ"),                        //
      //.SATA_EIDLE_VAL                 ( 3'b100),                              //
      //.SATA_MAX_BURST                 ( 8),                                   //
      //.SATA_MAX_INIT                  (21),                                   //
      //.SATA_MAX_WAKE                  ( 7),                                   //
      //.SATA_MIN_BURST                 ( 4),                                   //
      //.SATA_MIN_INIT                  (12),                                   //
      //.SATA_MIN_WAKE                  ( 4),                                   //  
                                                                                
        //---------- MISC ------------------------------------------------------               
        .DMONITOR_CFG                   (24'h000B01),                           // Optimized for debug
        .RX_DEBUG_CFG                   (12'd0)                                 // Optimized for GES
      //.TST_RSV                        (32'd0),                                //
      //.UCODEER_CLR                    ( 1'd0)                                 //
                                                                                
    )                                                                           
    model_ap2_tst_gtxe2_channel_i                                                                     
    (                                                                           
                                                                                
        //---------- Clock -----------------------------------------------------                
        .GTGREFCLK                      (1'd0),                                 //
        .GTREFCLK0                      (GT_GTREFCLK0),                         //
        .GTREFCLK1                      (1'd0),                                 //
        .GTNORTHREFCLK0                 (1'd0),                                 //
        .GTNORTHREFCLK1                 (1'd0),                                 //
        .GTSOUTHREFCLK0                 (1'd0),                                 //
        .GTSOUTHREFCLK1                 (1'd0),                                 //
        .QPLLCLK                        (GT_QPLLCLK),                           //
        .QPLLREFCLK                     (GT_QPLLREFCLK),                        //
        .TXUSRCLK                       (GT_TXUSRCLK),                          //
        .RXUSRCLK                       (GT_RXUSRCLK),                          //
        .TXUSRCLK2                      (GT_TXUSRCLK2),                         //
        .RXUSRCLK2                      (GT_RXUSRCLK2),                         //
        .TXSYSCLKSEL                    (GT_TXSYSCLKSEL),                       // 
        .RXSYSCLKSEL                    (GT_RXSYSCLKSEL),                       // 
        .TXOUTCLKSEL                    (txoutclksel),                          //
        .RXOUTCLKSEL                    (rxoutclksel),                          //
        .CPLLREFCLKSEL                  (3'd1),                                 //
        .CPLLLOCKDETCLK                 (1'd0),                                 //
        .CPLLLOCKEN                     (1'd1),                                 // 
        .CLKRSVD                        ({2'd0, dmonitorclk, GT_OOBCLK}),       // Optimized for debug
                                                                                
        .TXOUTCLK                       (GT_TXOUTCLK),                          //
        .RXOUTCLK                       (GT_RXOUTCLK),                          //
        .TXOUTCLKFABRIC                 (),                                     //
        .RXOUTCLKFABRIC                 (),                                     //
        .TXOUTCLKPCS                    (),                                     //
        .RXOUTCLKPCS                    (),                                     //
        .CPLLLOCK                       (GT_CPLLLOCK),                          //
        .CPLLREFCLKLOST                 (),                                     //
        .CPLLFBCLKLOST                  (),                                     //
        .RXCDRLOCK                      (GT_RXCDRLOCK),                         //
        .GTREFCLKMONITOR                (),                                     //
                                                                                
        //---------- Reset -----------------------------------------------------                
        .CPLLPD                         (cpllpd | GT_CPLLPD),                   // 
        .CPLLRESET                      (cpllrst | GT_CPLLRESET),               //
        .TXUSERRDY                      (GT_TXUSERRDY),                         //
        .RXUSERRDY                      (GT_RXUSERRDY),                         //
        .CFGRESET                       (1'd0),                                 //
        .GTRESETSEL                     (1'd0),                                 //
        .RESETOVRD                      (GT_RESETOVRD),                         //
        .GTTXRESET                      (GT_GTTXRESET),                         //
        .GTRXRESET                      (GT_GTRXRESET),                         //
                                                                               
        .TXRESETDONE                    (GT_TXRESETDONE),                       //
        .RXRESETDONE                    (GT_RXRESETDONE),                       //
                                                                                
        //---------- TX Data ---------------------------------------------------                
        .TXDATA                         ({32'd0, GT_TXDATA}),                   //
        .TXCHARISK                      ({ 4'd0, GT_TXDATAK}),                  //
                                                                                
        .GTXTXP                         (GT_TXP),                               // GTX
        .GTXTXN                         (GT_TXN),                               // GTX
                                                                                
        //---------- RX Data ---------------------------------------------------                
        .GTXRXP                         (GT_RXP),                               // GTX
        .GTXRXN                         (GT_RXN),                               // GTX
                                                                                
        .RXDATA                         (rxdata),                               //
        .RXCHARISK                      (rxdatak),                              //
                                                                                
        //---------- Command ---------------------------------------------------                
        .TXDETECTRX                     (GT_TXDETECTRX),                        //
        .TXPDELECIDLEMODE               ( 1'd0),                                //
        .RXELECIDLEMODE                 ( 2'd0),                                //
        .TXELECIDLE                     (GT_TXELECIDLE),                        //
        .TXCHARDISPMODE                 ({7'd0, GT_TXCOMPLIANCE}),              //
        .TXCHARDISPVAL                  ( 8'd0),                                //
        .TXPOLARITY                     ( 1'b0),                                //
        .RXPOLARITY                     (GT_RXPOLARITY),                        //
        .TXPD                           (GT_TXPOWERDOWN),                       //
        .RXPD                           (GT_RXPOWERDOWN),                       //
        .TXRATE                         (GT_TXRATE),                            //
        .RXRATE                         (GT_RXRATE),                            //
                                                                                
        //---------- Electrical Command ----------------------------------------                
        .TXMARGIN                       (GT_TXMARGIN),                          //
        .TXSWING                        (GT_TXSWING),                           //
        .TXDEEMPH                       (GT_TXDEEMPH),                          //
        .TXINHIBIT                      (1'd0),                                 // 
        .TXBUFDIFFCTRL                  (3'b100),                               // 
        .TXDIFFCTRL                     (4'b1100),                              //   
        .TXPRECURSOR                    (GT_TXPRECURSOR),                       // 
        .TXPRECURSORINV                 (1'd0),                                 // 
        .TXMAINCURSOR                   (GT_TXMAINCURSOR),                      // 
        .TXPOSTCURSOR                   (GT_TXPOSTCURSOR),                      // 
        .TXPOSTCURSORINV                (1'd0),                                 // 
                                                                                
        //---------- Status ----------------------------------------------------                
        .RXVALID                        (GT_RXVALID),                           //
        .PHYSTATUS                      (GT_PHYSTATUS),                         //
        .RXELECIDLE                     (GT_RXELECIDLE),                        // 
        .RXSTATUS                       (GT_RXSTATUS),                          //
        .TXRATEDONE                     (GT_TXRATEDONE),                        //
        .RXRATEDONE                     (GT_RXRATEDONE),                        //
                                                                                
        //---------- DRP -------------------------------------------------------                
        .DRPCLK                         (GT_DRPCLK),                            //
        .DRPADDR                        (GT_DRPADDR),                           //
        .DRPEN                          (GT_DRPEN),                             //
        .DRPDI                          (GT_DRPDI),                             //
        .DRPWE                          (GT_DRPWE),                             //
                                                                                
        .DRPDO                          (GT_DRPDO),                             //
        .DRPRDY                         (GT_DRPRDY),                            //
                                                                                
        //---------- PMA -------------------------------------------------------                
        .TXPMARESET                     (GT_TXPMARESET),                        //
        .RXPMARESET                     (GT_RXPMARESET),                        //
        .RXLPMEN                        (rxlpmen),                              // 
        .RXLPMHFHOLD                    ( 1'd0),                                // 
        .RXLPMHFOVRDEN                  ( 1'd0),                                // 
        .RXLPMLFHOLD                    ( 1'd0),                                // 
        .RXLPMLFKLOVRDEN                ( 1'd0),                                // 
        .TXQPIBIASEN                    ( 1'd0),                                // 
        .TXQPISTRONGPDOWN               ( 1'd0),                                // 
        .TXQPIWEAKPUP                   ( 1'd0),                                // 
        .RXQPIEN                        ( 1'd0),                                // 
        .PMARSVDIN                      ( 5'd0),                                // 
        .PMARSVDIN2                     ( 5'd0),                                // GTX 
        .GTRSVD                         (16'd0),                                // 
                                                                                
        .TXQPISENP                      (),                                     // 
        .TXQPISENN                      (),                                     // 
        .RXQPISENP                      (),                                     // 
        .RXQPISENN                      (),                                     // 
        .DMONITOROUT                    (dmonitorout[7:0]),                     // GTX 8-bits
                                                                                
        //---------- PCS -------------------------------------------------------                
        .TXPCSRESET                     (GT_TXPCSRESET),                        //
        .RXPCSRESET                     (GT_RXPCSRESET),                        //
        .PCSRSVDIN                      (16'd0),                                // [0]: 1 = TXRATE async, [1]: 1 = RXRATE async  
        .PCSRSVDIN2                     ( 5'd0),                                // 
                                                                                
        .PCSRSVDOUT                     (),                                     // 
        //---------- CDR -------------------------------------------------------                
        .RXCDRRESET                     (GT_RXCDRRESET),                        //
        .RXCDRRESETRSV                  (1'd0),                                 // 
        .RXCDRFREQRESET                 (GT_RXCDRFREQRESET),                    // 
        .RXCDRHOLD                      (1'b0),                                 //
        .RXCDROVRDEN                    (1'd0),                                 // 
                                                                                
        //---------- DFE -------------------------------------------------------                
        .RXDFELPMRESET                  (GT_RXDFELPMRESET),                     //  
        .RXDFECM1EN                     (1'd0),                                 // 
        .RXDFEVSEN                      (1'd0),                                 // 
        .RXDFETAP2HOLD                  (1'd0),                                 // 
        .RXDFETAP2OVRDEN                (1'd0),                                 // 
        .RXDFETAP3HOLD                  (1'd0),                                 // 
        .RXDFETAP3OVRDEN                (1'd0),                                 // 
        .RXDFETAP4HOLD                  (1'd0),                                 // 
        .RXDFETAP4OVRDEN                (1'd0),                                 // 
        .RXDFETAP5HOLD                  (1'd0),                                 // 
        .RXDFETAP5OVRDEN                (1'd0),                                 // 
        .RXDFEAGCHOLD                   (GT_RX_CONVERGE),                       // Optimized for GES, Set to 1 after convergence 
        .RXDFEAGCOVRDEN                 (1'd0),                                 // 
        .RXDFELFHOLD                    (1'd0),                                 // 
        .RXDFELFOVRDEN                  (1'd1),                                 // Optimized for GES
        .RXDFEUTHOLD                    (1'd0),                                 // 
        .RXDFEUTOVRDEN                  (1'd0),                                 // 
        .RXDFEVPHOLD                    (1'd0),                                 // 
        .RXDFEVPOVRDEN                  (1'd0),                                 // 
        .RXDFEXYDEN                     (1'd0),                                 // 
        .RXDFEXYDHOLD                   (1'd0),                                 // GTX 
        .RXDFEXYDOVRDEN                 (1'd0),                                 // GTX
        .RXMONITORSEL                   (2'd0),                                 //
                                                                                
        .RXMONITOROUT                   (),                                     // 
             
        //---------- OS --------------------------------------------------------         
        .RXOSHOLD                       (1'd0),                                 // 
        .RXOSOVRDEN                     (1'd0),                                 //        
                                                                                
        //---------- Eye Scan --------------------------------------------------                
        .EYESCANRESET                   (GT_EYESCANRESET),                      // 
        .EYESCANMODE                    (1'd0),                                 // 
        .EYESCANTRIGGER                 (1'b0),                                 //
                                                                                
        .EYESCANDATAERROR               (GT_EYESCANDATAERROR),                  //
                                                                                
        //---------- TX Buffer -------------------------------------------------                
        .TXBUFSTATUS                    (),                                     //
                                                                                
        //---------- RX Buffer -------------------------------------------------                
        .RXBUFRESET                     (GT_RXBUFRESET),                        //
                                                                                
        .RXBUFSTATUS                    (GT_RXBUFSTATUS),                       //
                                                                                
        //---------- TX Sync ---------------------------------------------------                
        .TXPHDLYRESET                   (1'd0),                                 //
        .TXPHDLYTSTCLK                  (1'd0),                                 //
        .TXPHALIGN                      (GT_TXPHALIGN),                         // 
        .TXPHALIGNEN                    (GT_TXPHALIGNEN),                       //  
        .TXPHDLYPD                      (1'd0),                                 // 
        .TXPHINIT                       (GT_TXPHINIT),                          //  
        .TXPHOVRDEN                     (1'd0),                                 //
        .TXDLYBYPASS                    (GT_TXDLYBYPASS),                       //  
        .TXDLYSRESET                    (GT_TXDLYSRESET),                       // 
        .TXDLYEN                        (GT_TXDLYEN),                           //  
        .TXDLYOVRDEN                    (1'd0),                                 //
        .TXDLYHOLD                      (1'd0),                                 // 
        .TXDLYUPDOWN                    (1'd0),                                 //
                                                                                
        .TXPHALIGNDONE                  (GT_TXPHALIGNDONE),                     // 
        .TXPHINITDONE                   (GT_TXPHINITDONE),                      // 
        .TXDLYSRESETDONE                (GT_TXDLYSRESETDONE),                   //
                                                                                
        //---------- RX Sync ---------------------------------------------------                  
        .RXPHDLYRESET                   (1'd0),                                 //
        .RXPHALIGN                      (GT_RXPHALIGN),                         //
        .RXPHALIGNEN                    (GT_RXPHALIGNEN),                       //
        .RXPHDLYPD                      (1'd0),                                 // 
        .RXPHOVRDEN                     (1'd0),                                 // 
        .RXDLYBYPASS                    (GT_RXDLYBYPASS),                       //  
        .RXDLYSRESET                    (GT_RXDLYSRESET),                       // 
        .RXDLYEN                        (GT_RXDLYEN),                           // 
        .RXDLYOVRDEN                    (1'd0),                                 //
        .RXDDIEN                        (GT_RXDDIEN),                           //
                                                                                
        .RXPHALIGNDONE                  (GT_RXPHALIGNDONE),                     //  
        .RXPHMONITOR                    (),                                     //
        .RXPHSLIPMONITOR                (),                                     // 
        .RXDLYSRESETDONE                (GT_RXDLYSRESETDONE),                   // 
                                                                                
        //---------- Comma Alignment -------------------------------------------                 
        .RXCOMMADETEN                   ( 1'd1),                                //
        .RXMCOMMAALIGNEN                (!GT_GEN3),                             // 0 = disable comma alignment in Gen3
        .RXPCOMMAALIGNEN                (!GT_GEN3),                             // 0 = disable comma alignment in Gen3
        .RXSLIDE                        ( GT_RXSLIDE),                          //
                                                                                
        .RXCOMMADET                     (GT_RXCOMMADET),                        //
        .RXCHARISCOMMA                  (rxchariscomma),                        // 
        .RXBYTEISALIGNED                (GT_RXBYTEISALIGNED),                   //
        .RXBYTEREALIGN                  (GT_RXBYTEREALIGN),                     //
                                                                                
        //---------- Channel Bonding -------------------------------------------                
        .RXCHBONDEN                     (GT_RXCHBONDEN),                        //
        .RXCHBONDI                      (GT_RXCHBONDI),                         //
        .RXCHBONDLEVEL                  (GT_RXCHBONDLEVEL),                     //
        .RXCHBONDMASTER                 (GT_RXCHBONDMASTER),                    //
        .RXCHBONDSLAVE                  (GT_RXCHBONDSLAVE),                     //
                                                                                
        .RXCHANBONDSEQ                  (),                                     //
        .RXCHANISALIGNED                (GT_RXCHANISALIGNED),                   //
        .RXCHANREALIGN                  (),                                     //
        .RXCHBONDO                      (GT_RXCHBONDO),                         //
                                                                                
        //---------- Clock Correction  -----------------------------------------                
        .RXCLKCORCNT                    (),                                     //
                                                                                
        //---------- 8b10b -----------------------------------------------------                
        .TX8B10BBYPASS                  (8'd0),                                 //
        .TX8B10BEN                      (!GT_GEN3),                             // 0 = disable TX 8b10b in Gen3
        .RX8B10BEN                      (!GT_GEN3),                             // 0 = disable RX 8b10b in Gen3
                                                                                
        .RXDISPERR                      (GT_RXDISPERR),                         //
        .RXNOTINTABLE                   (GT_RXNOTINTABLE),                      //
                                                                                
        //---------- 64b/66b & 64b/67b -----------------------------------------                  
        .TXHEADER                       (3'd0),                                 //
        .TXSEQUENCE                     (7'd0),                                 //
        .TXSTARTSEQ                     (1'd0),                                 //                                                              
        .RXGEARBOXSLIP                  (1'd0),                                 //
                                                                                
        .TXGEARBOXREADY                 (),                                     // 
        .RXDATAVALID                    (),                                     //
        .RXHEADER                       (),                                     //
        .RXHEADERVALID                  (),                                     //
        .RXSTARTOFSEQ                   (),                                     //
                                                                                
        //---------- PRBS/Loopback ---------------------------------------------                
        .TXPRBSSEL                      (GT_TXPRBSSEL),                         //
        .RXPRBSSEL                      (GT_RXPRBSSEL),                         //
        .TXPRBSFORCEERR                 (GT_TXPRBSFORCEERR),                    //
        .RXPRBSCNTRESET                 (GT_RXPRBSCNTRESET),                    // 
        .LOOPBACK                       (GT_LOOPBACK),                          // 
                                                                                
        .RXPRBSERR                      (GT_RXPRBSERR),                         //
                                                                                
        //---------- OOB -------------------------------------------------------                
        .TXCOMINIT                      (1'd0),                                 //
        .TXCOMSAS                       (1'd0),                                 //
        .TXCOMWAKE                      (1'd0),                                 //
        .RXOOBRESET                     (1'd0),                                 // 
                                                                                
        .TXCOMFINISH                    (),                                     //
        .RXCOMINITDET                   (),                                     //
        .RXCOMSASDET                    (),                                     //
        .RXCOMWAKEDET                   (),                                     //
                                                                                
        //---------- MISC ------------------------------------------------------                
        .SETERRSTATUS                   ( 1'd0),                                // 
        .TXDIFFPD                       ( 1'd0),                                // 
        .TXPISOPD                       ( 1'd0),                                // 
        .TSTIN                          (20'hFFFFF),                            //  
                                                                                
        .TSTOUT                         ()                                      // GTX
    
    );
    
    //---------- Default -------------------------------------------------------
    assign dmonitorout[14:8] = 7'd0;                                            // GTH GTP
    assign GT_TXSYNCOUT      = 1'd0;                                            // GTH GTP  
    assign GT_TXSYNCDONE     = 1'd0;                                            // GTH GTP 
    assign GT_RXSYNCOUT      = 1'd0;                                            // GTH GTP
    assign GT_RXSYNCDONE     = 1'd0;                                            // GTH GTP
    assign GT_RXPMARESETDONE = 1'd0;                                            // GTH GTP               
            
    end

endgenerate
    
//---------- GT Wrapper Outputs ------------------------------------------------
assign GT_RXDATA        = rxdata [31:0];
assign GT_RXDATAK       = rxdatak[ 3:0];
assign GT_RXCHARISCOMMA = rxchariscomma[ 3:0];
assign GT_DMONITOROUT   = dmonitorout;

endmodule



`timescale 1ns/1ps
module model_ap2_tst_gtx_cpllpd_ovrd (                                                                                        
    input   i_ibufds_gte2,                                                                                     
    output  o_cpllpd_ovrd,                                                                                     
    output  o_cpllreset_ovrd                                                                                   
    );                                                                                                         
    (* equivalent_register_removal="no" *)  reg [95:0] cpllpd_wait = 96'hFFFFFFFFFFFFFFFFFFFFFFFF;             
    (* equivalent_register_removal="no" *)  reg [127:0] cpllreset_wait = 128'h000000000000000000000000000000FF;
    always @(posedge i_ibufds_gte2)                                                                            
    begin                                                                                                      
        cpllpd_wait <= {cpllpd_wait[94:0], 1'b0};                                                              
        cpllreset_wait <= {cpllreset_wait[126:0], 1'b0};                                                       
    end                                                                                                        
    assign o_cpllpd_ovrd = cpllpd_wait[95];                                                                    
    assign o_cpllreset_ovrd = cpllreset_wait[127];                                                             
endmodule


module model_ap2_tst_pipe_clock #
(

    parameter PCIE_ASYNC_EN      = "FALSE",                 // PCIe async enable
    parameter PCIE_TXBUF_EN      = "FALSE",                 // PCIe TX buffer enable for Gen1/Gen2 only
    parameter PCIE_CLK_SHARING_EN= "FALSE",                 // Enable Clock Sharing
    parameter PCIE_LANE          = 1,                       // PCIe number of lanes
    parameter PCIE_LINK_SPEED    = 3,                       // PCIe link speed 
    parameter PCIE_REFCLK_FREQ   = 0,                       // PCIe reference clock frequency
    parameter PCIE_USERCLK1_FREQ = 2,                       // PCIe user clock 1 frequency
    parameter PCIE_USERCLK2_FREQ = 2,                       // PCIe user clock 2 frequency
    parameter PCIE_OOBCLK_MODE   = 1,                       // PCIe oob clock mode
    parameter PCIE_DEBUG_MODE    = 0                        // PCIe Debug mode
    
)

(

    //---------- Input -------------------------------------
    input                       CLK_CLK,
    input                       CLK_TXOUTCLK,
    input       [PCIE_LANE-1:0] CLK_RXOUTCLK_IN,
    input                       CLK_RST_N,
    input       [PCIE_LANE-1:0] CLK_PCLK_SEL,
    input       [PCIE_LANE-1:0] CLK_PCLK_SEL_SLAVE,
    input                       CLK_GEN3,
    
    //---------- Output ------------------------------------
    output                      CLK_PCLK,
    output                      CLK_PCLK_SLAVE,
    output                      CLK_RXUSRCLK,
    output      [PCIE_LANE-1:0] CLK_RXOUTCLK_OUT,
    output                      CLK_DCLK,
    output                      CLK_OOBCLK,
    output                      CLK_USERCLK1,
    output                      CLK_USERCLK2,
    output                      CLK_MMCM_LOCK
    
);
    
    //---------- Select Clock Divider ----------------------
    localparam          DIVCLK_DIVIDE    = (PCIE_REFCLK_FREQ == 2) ? 1 :
                                           (PCIE_REFCLK_FREQ == 1) ? 1 : 1;
                                               
    localparam          CLKFBOUT_MULT_F  = (PCIE_REFCLK_FREQ == 2) ? 4 :
                                           (PCIE_REFCLK_FREQ == 1) ? 8 : 10;
               
    localparam          CLKIN1_PERIOD    = (PCIE_REFCLK_FREQ == 2) ? 4 :
                                           (PCIE_REFCLK_FREQ == 1) ? 8 : 10;
                                               
    localparam          CLKOUT0_DIVIDE_F = 8;
    
    localparam          CLKOUT1_DIVIDE   = 4;
    
    localparam          CLKOUT2_DIVIDE   = (PCIE_USERCLK1_FREQ == 5) ?  2 : 
                                           (PCIE_USERCLK1_FREQ == 4) ?  4 :
                                           (PCIE_USERCLK1_FREQ == 3) ?  8 :
                                           (PCIE_USERCLK1_FREQ == 1) ? 32 : 16;
                                               
    localparam          CLKOUT3_DIVIDE   = (PCIE_USERCLK2_FREQ == 5) ?  2 : 
                                           (PCIE_USERCLK2_FREQ == 4) ?  4 :
                                           (PCIE_USERCLK2_FREQ == 3) ?  8 :
                                           (PCIE_USERCLK2_FREQ == 1) ? 32 : 16;
                                           
    localparam          CLKOUT4_DIVIDE   = 20;

    localparam          PCIE_GEN1_MODE    = 1'b0;             // PCIe link speed is GEN1 only
                                    
       
    //---------- Input Registers ---------------------------
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0] pclk_sel_reg1 = {PCIE_LANE{1'd0}};
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0] pclk_sel_slave_reg1 = {PCIE_LANE{1'd0}};
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                         gen3_reg1     = 1'd0;
    
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0] pclk_sel_reg2 = {PCIE_LANE{1'd0}};
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg         [PCIE_LANE-1:0] pclk_sel_slave_reg2 = {PCIE_LANE{1'd0}};
(* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *)    reg                         gen3_reg2     = 1'd0;   
       
    //---------- Internal Signals -------------------------- 
    wire                            refclk;
    wire                            mmcm_fb;
    wire                            clk_125mhz;
    wire                            clk_125mhz_buf;
    wire                            clk_250mhz;
    wire                            userclk1;
    wire                            userclk2;
    wire                            oobclk;
    reg    pclk_sel = 1'd0;
    reg                             pclk_sel_slave = 1'd0;

    //---------- Output Registers --------------------------
    wire                        pclk_1;
    wire                        pclk;
    wire                        userclk1_1;
    wire                        userclk2_1;
    wire                        mmcm_lock;
    
    //---------- Generate Per-Lane Signals -----------------
    genvar              i;                                  // Index for per-lane signals



//---------- Input FF ----------------------------------------------------------
always @ (posedge pclk)
begin

    if (!CLK_RST_N)
        begin
        //---------- 1st Stage FF --------------------------
        pclk_sel_reg1 <= {PCIE_LANE{1'd0}};
        pclk_sel_slave_reg1 <= {PCIE_LANE{1'd0}};
        gen3_reg1     <= 1'd0;
        //---------- 2nd Stage FF --------------------------
        pclk_sel_reg2 <= {PCIE_LANE{1'd0}};
        pclk_sel_slave_reg2 <= {PCIE_LANE{1'd0}};
        gen3_reg2     <= 1'd0;
        end
    else
        begin  
        //---------- 1st Stage FF --------------------------
        pclk_sel_reg1 <= CLK_PCLK_SEL;
        pclk_sel_slave_reg1 <= CLK_PCLK_SEL_SLAVE;
        gen3_reg1     <= CLK_GEN3;
        //---------- 2nd Stage FF --------------------------
        pclk_sel_reg2 <= pclk_sel_reg1;
        pclk_sel_slave_reg2 <= pclk_sel_slave_reg1;
        gen3_reg2     <= gen3_reg1;
        end
        
end


   
//---------- Select Reference clock or TXOUTCLK --------------------------------   
generate if ((PCIE_TXBUF_EN == "TRUE") && (PCIE_LINK_SPEED != 3))

    begin : refclk_i

    //---------- Select Reference Clock ----------------------------------------
    BUFG refclk_i
    (
    
        //---------- Input -------------------------------------
        .I                          (CLK_CLK),
        //---------- Output ------------------------------------
        .O                          (refclk)
       
    );
      
    end

else

    begin : txoutclk_i
    
    //---------- Select TXOUTCLK -----------------------------------------------
    BUFG txoutclk_i
    (
    
        //---------- Input -------------------------------------
        .I                          (CLK_TXOUTCLK),
        //---------- Output ------------------------------------
        .O                          (refclk)
       
    );
   
    end

endgenerate



//---------- MMCM --------------------------------------------------------------
MMCME2_ADV #
(

    .BANDWIDTH                  ("OPTIMIZED"),
    .CLKOUT4_CASCADE            ("FALSE"),
    .COMPENSATION               ("ZHOLD"),
    .STARTUP_WAIT               ("FALSE"),
    .DIVCLK_DIVIDE              (DIVCLK_DIVIDE),
    .CLKFBOUT_MULT_F            (CLKFBOUT_MULT_F),  
    .CLKFBOUT_PHASE             (0.000),
    .CLKFBOUT_USE_FINE_PS       ("FALSE"),
    .CLKOUT0_DIVIDE_F           (CLKOUT0_DIVIDE_F),                    
    .CLKOUT0_PHASE              (0.000),
    .CLKOUT0_DUTY_CYCLE         (0.500),
    .CLKOUT0_USE_FINE_PS        ("FALSE"),
    .CLKOUT1_DIVIDE             (CLKOUT1_DIVIDE),                    
    .CLKOUT1_PHASE              (0.000),
    .CLKOUT1_DUTY_CYCLE         (0.500),
    .CLKOUT1_USE_FINE_PS        ("FALSE"),
    .CLKOUT2_DIVIDE             (CLKOUT2_DIVIDE),                  
    .CLKOUT2_PHASE              (0.000),
    .CLKOUT2_DUTY_CYCLE         (0.500),
    .CLKOUT2_USE_FINE_PS        ("FALSE"),
    .CLKOUT3_DIVIDE             (CLKOUT3_DIVIDE),                  
    .CLKOUT3_PHASE              (0.000),
    .CLKOUT3_DUTY_CYCLE         (0.500),
    .CLKOUT3_USE_FINE_PS        ("FALSE"),
    .CLKOUT4_DIVIDE             (CLKOUT4_DIVIDE),                  
    .CLKOUT4_PHASE              (0.000),
    .CLKOUT4_DUTY_CYCLE         (0.500),
    .CLKOUT4_USE_FINE_PS        ("FALSE"),
    .CLKIN1_PERIOD              (CLKIN1_PERIOD),                   
    .REF_JITTER1                (0.010)
    
)
mmcm_i
(

     //---------- Input ------------------------------------
    .CLKIN1                     (refclk),
    .CLKIN2                     (1'd0),                     // not used, comment out CLKIN2 if it cause implementation issues
  //.CLKIN2                     (refclk),                   // not used, comment out CLKIN2 if it cause implementation issues
    .CLKINSEL                   (1'd1),
    .CLKFBIN                    (mmcm_fb),
    .RST                        (!CLK_RST_N),
    .PWRDWN                     (1'd0), 
    
    //---------- Output ------------------------------------
    .CLKFBOUT                   (mmcm_fb),
    .CLKFBOUTB                  (),
    .CLKOUT0                    (clk_125mhz),
    .CLKOUT0B                   (),
    .CLKOUT1                    (clk_250mhz),
    .CLKOUT1B                   (),
    .CLKOUT2                    (userclk1),
    .CLKOUT2B                   (),
    .CLKOUT3                    (userclk2),
    .CLKOUT3B                   (),
    .CLKOUT4                    (oobclk),
    .CLKOUT5                    (),
    .CLKOUT6                    (),
    .LOCKED                     (mmcm_lock),
    
    //---------- Dynamic Reconfiguration -------------------
    .DCLK                       ( 1'd0),
    .DADDR                      ( 7'd0),
    .DEN                        ( 1'd0),
    .DWE                        ( 1'd0),
    .DI                         (16'd0),
    .DO                         (),
    .DRDY                       (),
    
    //---------- Dynamic Phase Shift -----------------------
    .PSCLK                      (1'd0),
    .PSEN                       (1'd0),
    .PSINCDEC                   (1'd0),
    .PSDONE                     (),
    
    //---------- Status ------------------------------------
    .CLKINSTOPPED               (),
    .CLKFBSTOPPED               ()  

); 
  


//---------- Select PCLK MUX ---------------------------------------------------
generate if (PCIE_LINK_SPEED != 1) 

    begin : pclk_i1_bufgctrl
    //---------- PCLK Mux ----------------------------------
    BUFGCTRL pclk_i1
    (
        //---------- Input ---------------------------------
        .CE0                        (1'd1),         
        .CE1                        (1'd1),        
        .I0                         (clk_125mhz),   
        .I1                         (clk_250mhz),   
        .IGNORE0                    (1'd0),        
        .IGNORE1                    (1'd0),        
        .S0                         (~pclk_sel),    
        .S1                         ( pclk_sel),    
        //---------- Output --------------------------------
        .O                          (pclk_1)
    );
    end

else 

    //---------- Select PCLK Buffer ------------------------
    begin : pclk_i1_bufg
    //---------- PCLK Buffer -------------------------------
    BUFG pclk_i1
    (
        //---------- Input ---------------------------------
        .I                          (clk_125mhz), 
        //---------- Output --------------------------------
        .O                          (clk_125mhz_buf)
    );
    assign pclk_1 = clk_125mhz_buf;
    end 

endgenerate

//---------- Select PCLK MUX for Slave---------------------------------------------------
generate  if(PCIE_CLK_SHARING_EN == "FALSE")
   //---------- PCLK MUX for Slave------------------// 
    begin : pclk_slave_disable
    assign CLK_PCLK_SLAVE = 1'b0;
    end  

else if (PCIE_LINK_SPEED != 1) 

    begin : pclk_slave_bufgctrl
    //---------- PCLK Mux ----------------------------------
    BUFGCTRL pclk_slave
    (
        //---------- Input ---------------------------------
        .CE0                        (1'd1),         
        .CE1                        (1'd1),        
        .I0                         (clk_125mhz),   
        .I1                         (clk_250mhz),   
        .IGNORE0                    (1'd0),        
        .IGNORE1                    (1'd0),        
        .S0                         (~pclk_sel_slave),    
        .S1                         ( pclk_sel_slave),    
        //---------- Output --------------------------------
        .O                          (CLK_PCLK_SLAVE)
    );
    end

else 

    //---------- Select PCLK Buffer ------------------------
    begin : pclk_slave_bufg
    //---------- PCLK Buffer -------------------------------
    BUFG pclk_slave
    (
        //---------- Input ---------------------------------
        .I                          (clk_125mhz), 
        //---------- Output --------------------------------
        .O                          (CLK_PCLK_SLAVE)
    );
    end 

endgenerate



//---------- Generate RXOUTCLK Buffer for Debug --------------------------------
generate if ((PCIE_DEBUG_MODE == 1) || (PCIE_ASYNC_EN == "TRUE"))
        
    begin : rxoutclk_per_lane
    //---------- Generate per Lane -------------------------
    for (i=0; i<PCIE_LANE; i=i+1) 
    
        begin : rxoutclk_i
        //---------- RXOUTCLK Buffer -----------------------
        BUFG rxoutclk_i
        (
            //---------- Input -----------------------------
            .I                          (CLK_RXOUTCLK_IN[i]), 
            //---------- Output ----------------------------
            .O                          (CLK_RXOUTCLK_OUT[i])
        );
        end

    end 
        
else

    //---------- Disable RXOUTCLK Buffer for Normal Operation 
    begin : rxoutclk_i_disable
    assign CLK_RXOUTCLK_OUT = {PCIE_LANE{1'd0}};
    end       
            
endgenerate 


//---------- Generate DCLK Buffer ----------------------------------------------
//generate if (PCIE_USERCLK2_FREQ <= 3)
//---------- Disable DCLK Buffer -----------------------
//    begin : dclk_i
//    assign CLK_DCLK = userclk2_1;                       // always less than 125Mhz
//   end
//else
//    begin : dclk_i_bufg
//---------- DCLK Buffer -------------------------------
//    BUFG dclk_i
//    (
//---------- Input ---------------------------------
//        .I                          (clk_125mhz), 
//---------- Output --------------------------------
//        .O                          (CLK_DCLK)
//    );
//    end 
//endgenerate

generate if (PCIE_LINK_SPEED != 1)

    begin : dclk_i_bufg
    //---------- DCLK Buffer -------------------------------
    BUFG dclk_i
    (
        //---------- Input ---------------------------------
        .I                          (clk_125mhz),
        //---------- Output --------------------------------
        .O                          (CLK_DCLK)
    );
    end

else

    //---------- Disable DCLK Buffer -----------------------
    begin : dclk_i
    assign CLK_DCLK = clk_125mhz_buf;                       // always 125 MHz in Gen1
    end

endgenerate




//---------- Generate USERCLK1 Buffer ------------------------------------------
generate if (PCIE_GEN1_MODE == 1'b1 && PCIE_USERCLK1_FREQ == 3) 
    //---------- USERCLK1 same as PCLK -------------------
    begin :userclk1_i1_no_bufg
    assign userclk1_1 = pclk_1;
    end 
else
    begin : userclk1_i1
    //---------- USERCLK1 Buffer ---------------------------
    BUFG usrclk1_i1
    (
        //---------- Input ---------------------------------
        .I                          (userclk1),
        //---------- Output --------------------------------
        .O                          (userclk1_1)
    );
    end 
endgenerate 



//---------- Generate USERCLK2 Buffer ------------------------------------------

generate if (PCIE_GEN1_MODE == 1'b1 && PCIE_USERCLK2_FREQ == 3 ) 
//---------- USERCLK2 same as PCLK -------------------
    begin : userclk2_i1_no_bufg0
    assign userclk2_1 = pclk_1;
    end 
else if (PCIE_USERCLK2_FREQ == PCIE_USERCLK1_FREQ ) 
//---------- USERCLK2 same as USERCLK1 -------------------
    begin : userclk2_i1_no_bufg1
    assign userclk2_1 = userclk1_1;
    end  
else    
    begin : userclk2_i1
    //---------- USERCLK2 Buffer ---------------------------
    BUFG usrclk2_i1
    (
        //---------- Input ---------------------------------
        .I                          (userclk2),
        //---------- Output --------------------------------
        .O                          (userclk2_1)
    );
    end
endgenerate 



//---------- Generate OOBCLK Buffer --------------------------------------------
generate if (PCIE_OOBCLK_MODE == 2) 

    begin : oobclk_i1
    //---------- OOBCLK Buffer -----------------------------
    BUFG oobclk_i1
    (
        //---------- Input ---------------------------------
        .I                          (oobclk),
        //---------- Output --------------------------------
        .O                          (CLK_OOBCLK)
    );
    end

else 
        
    //---------- Disable OOBCLK Buffer ---------------------
    begin : oobclk_i1_disable
    assign CLK_OOBCLK = pclk;
    end  

endgenerate 


// Disabled Second Stage Buffers
    assign pclk         = pclk_1;
    assign CLK_RXUSRCLK = pclk_1;
    assign CLK_USERCLK1 = userclk1_1;
    assign CLK_USERCLK2 = userclk2_1;
 



//---------- Select PCLK -------------------------------------------------------
always @ (posedge pclk)
begin

    if (!CLK_RST_N)
        pclk_sel <= 1'd0;
    else
        begin 
        //---------- Select 250 MHz ------------------------
        if (&pclk_sel_reg2)
            pclk_sel <= 1'd1;
        //---------- Select 125 MHz ------------------------  
        else if (&(~pclk_sel_reg2))
            pclk_sel <= 1'd0;  
        //---------- Hold PCLK -----------------------------
        else
            pclk_sel <= pclk_sel;
        end

end        

always @ (posedge pclk)
begin

    if (!CLK_RST_N)
        pclk_sel_slave<= 1'd0;
    else
        begin 
        //---------- Select 250 MHz ------------------------
        if (&pclk_sel_slave_reg2)
            pclk_sel_slave <= 1'd1;
        //---------- Select 125 MHz ------------------------  
        else if (&(~pclk_sel_slave_reg2))
            pclk_sel_slave <= 1'd0;  
        //---------- Hold PCLK -----------------------------
        else
            pclk_sel_slave <= pclk_sel_slave;
        end

end     



//---------- PIPE Clock Output -------------------------------------------------
assign CLK_PCLK      = pclk;
assign CLK_MMCM_LOCK = mmcm_lock;



endmodule


//-----------------------------------------------------------------------------
// Project    : AXI Memory Mapped Bridge to PCI Express
// File       : BRAM_SDP_MACRO_model.v
// Version    : 2.8
//-----------------------------------------------------------------------------

module BRAM_SDP_MACRO_model (DO, 
                   DI, RDADDR, RDCLK, RDEN, REGCE, RST, WE, WRADDR, WRCLK, WREN); 

   parameter BRAM_SIZE = "18Kb"; 
   parameter DEVICE = "VIRTEX5";
   parameter DO_REG = 0;
   parameter INIT = 72'h0;
   parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
   parameter INIT_FILE = "NONE";
   parameter READ_WIDTH = 36;
   parameter SIM_COLLISION_CHECK = "ALL";
   parameter SIM_MODE = "SAFE"; // This parameter is valid only for Virtex5
   parameter SRVAL = 72'h0;
   parameter WRITE_MODE = "WRITE_FIRST";
   parameter WRITE_WIDTH = 36;


   localparam READ_P = ( (READ_WIDTH == 9) ||  (READ_WIDTH == 17) || (READ_WIDTH == 18) || (READ_WIDTH == 33) || (READ_WIDTH == 34) || (READ_WIDTH == 35) || (READ_WIDTH == 36) || (READ_WIDTH == 65) || (READ_WIDTH == 66) || (READ_WIDTH == 67) || (READ_WIDTH == 68) || (READ_WIDTH == 69) || (READ_WIDTH == 70) || (READ_WIDTH == 71) || (READ_WIDTH == 72) ) ? "TRUE" : "FALSE" ;
   localparam WRITE_P = ( (WRITE_WIDTH == 9) ||  (WRITE_WIDTH == 17) || (WRITE_WIDTH == 18) || (WRITE_WIDTH == 33) || (WRITE_WIDTH == 34) || (WRITE_WIDTH == 35) || (WRITE_WIDTH == 36) || (WRITE_WIDTH == 65) || (WRITE_WIDTH == 66) || (WRITE_WIDTH == 67) || (WRITE_WIDTH == 68) || (WRITE_WIDTH == 69) || (WRITE_WIDTH == 70) || (WRITE_WIDTH == 71) || (WRITE_WIDTH == 72) ) ? "TRUE" : "FALSE" ;

   localparam valid_width = ( (READ_WIDTH == 1 || READ_WIDTH == 2 || READ_WIDTH == 4 || READ_WIDTH == 8 || READ_WIDTH == 9 || READ_WIDTH == 16 || READ_WIDTH == 18 || READ_WIDTH == 32 || READ_WIDTH == 36 || READ_WIDTH == 64 || READ_WIDTH == 72) && (WRITE_WIDTH == 1 || WRITE_WIDTH == 2 || WRITE_WIDTH == 4 || WRITE_WIDTH == 8 || WRITE_WIDTH == 9 || WRITE_WIDTH == 16 || WRITE_WIDTH == 18 || WRITE_WIDTH == 32 || WRITE_WIDTH == 36 || WRITE_WIDTH == 64 || WRITE_WIDTH == 72)) ? "TRUE" : "FALSE";

   // Parameter Checks for invalid combinations
   initial 
   begin
     if (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6");
     else
       begin 
       $display("Attribute Syntax Error : The attribute DEVICE on BRAM_SDP_MACRO instance %m is set to %s.  Allowed values of this attribute are VIRTEX5, VIRTEX6, 7SERIES, SPARTAN6.", DEVICE);
       #1 $finish;
       end
     if( (DEVICE == "VIRTEX5") && (READ_WIDTH != WRITE_WIDTH)) 
       begin
       $display("Attribute Syntax Error : The attributes READ_WIDTH, WRITE_WIDTH on BRAM_SDP_MACRO instance %m are set to %d, %d.  To use BRAM_SDP_MACRO, READ_WIDTH must be equal to WRITE_WIDTH", READ_WIDTH, WRITE_WIDTH);
        #1 $finish;
       end
     if( (DEVICE == "VIRTEX6" || DEVICE == "SPARTAN6" || DEVICE == "7SERIES") && ((READ_WIDTH != WRITE_WIDTH) && (READ_WIDTH/WRITE_WIDTH !=2) && (WRITE_WIDTH/READ_WIDTH !=2) && (valid_width == "FALSE") ) ) 
       begin
       $display("Attribute Syntax Error : The attributes READ_WIDTH, WRITE_WIDTH on BRAM_SDP_MACRO instance %m are set to %d, %d.  To use BRAM_SDP_MACRO, one of the following conditions must be true-\n 1. READ_WIDTH must be equal to WRITE_WIDTH \n 2. If assymetric, READ_WIDTH and WRITE_WIDTH must have a ratio of 2.\n 3. If assymetric, READ_WIDTH and WRITE_WIDTH should have values 1, 2, 4, 8, 9, 16, 18, 32, 36, 64, 72.", READ_WIDTH, WRITE_WIDTH);
        #1 $finish;
       end
     if (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES")
     begin
       case ({WRITE_P, READ_P})

             {"FALSE", "TRUE"}: 
                begin 
                  $display("Port Width Mismatch on READ_WIDTH : The width READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  The parity bit(s) have not been written and hence cannot be read. ", READ_WIDTH);
                end
             {"TRUE", "FALSE"}: 
                begin 
                  $display("Port Width Mismatch on WRITE_WIDTH: The width WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  The parity bit(s) cannot be read ", WRITE_WIDTH);
	        end
       endcase
       if(BRAM_SIZE == "18Kb" || BRAM_SIZE == "36Kb") ;
       else
         begin
          $display("Attribute Syntax Error : The attribute BRAM_SIZE on BRAM_SDP_MACRO instance %m is set to %s.  Legal values for this attribute are 18Kb or 36Kb", BRAM_SIZE);
          #1 $finish;
       end
      if (READ_WIDTH == 0)
        begin 
          $display("Attribute Syntax Error : The attribute READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  This attribute must atleast be equal to 1.", READ_WIDTH);
           #1 $finish;
        end
      if ( READ_WIDTH > 36 && BRAM_SIZE == "18Kb" )
        begin 
          $display("Attribute Syntax Error : The attribute READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  For BRAM_SIZE of 18Kb, allowed values of this attribute are 1 to 36.", READ_WIDTH);
          #1 $finish;
        end
      if (READ_WIDTH > 72)
        begin 
          $display("Attribute Syntax Error : The attribute READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  Allowed values of this attribute are 1 to 36 for BRAM_SIZE of 18Kb and 1 to 72 for BRAM_SIZE of 36Kb.", READ_WIDTH);
          #1 $finish;
        end
      if (WRITE_WIDTH == 0)
        begin 
          $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  This attribute must atleast be equal to 1.", WRITE_WIDTH);
           #1 $finish;
        end
      if (WRITE_WIDTH > 36 && BRAM_SIZE == "18Kb" )
        begin 
          $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  For BRAM_SIZE of 18Kb, allowed values of this attribute are 1 to 36.", WRITE_WIDTH);
          #1 $finish;
        end
      if (WRITE_WIDTH > 72)
        begin 
           $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  Allowed values of this attribute are 1 to 36 for BRAM_SIZE of 18Kb and 1 to 72 for BRAM_SIZE of 36Kb.", WRITE_WIDTH);
           #1 $finish;
        end
     end // end checks Virtex5
     if (DEVICE == "SPARTAN6")
       begin
         if(BRAM_SIZE == "9Kb" || BRAM_SIZE == "18Kb") ;
         else
         begin
           $display("Attribute Syntax Error : The attribute BRAM_SIZE on BRAM_SDP_MACRO instance %m is set to %s.  Legal values for this attribute are 9Kb or 18Kb", BRAM_SIZE);
           #1 $finish;
         end
         if (READ_WIDTH == 0)
           begin 
             $display("Attribute Syntax Error : The attribute READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  This attribute must atleast be equal to 1.", READ_WIDTH);
             #1 $finish;
           end
         if (READ_WIDTH > 36)
           begin 
             $display("Attribute Syntax Error : The attribute READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  Allowed values of this attribute are 1 to 36 for BRAM_SIZE of 9Kb and 1 to 36 for BRAM_SIZE of 18Kb.", READ_WIDTH);
             #1 $finish;
           end
         if (WRITE_WIDTH == 0)
           begin 
             $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  This attribute must atleast be equal to 1.", WRITE_WIDTH);
             #1 $finish;
           end
         if (WRITE_WIDTH > 36)
           begin 
             $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  Allowed values of this attribute are 1 to 36 for BRAM_SIZE of 9Kb and 1 to 36 for BRAM_SIZE of 18Kb.", WRITE_WIDTH);
             #1 $finish;
           end
         if (((WRITE_WIDTH > 18 ||  READ_WIDTH > 18)  && (WRITE_WIDTH != READ_WIDTH)) && (BRAM_SIZE == "9Kb"))
           begin 
             $display("Attribute Syntax Error : The attribute WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d and the READ_WIDTH is set to %d.  For read or write widths greater than 18, the same port width must be used for read and write when in 9Kb mode.", WRITE_WIDTH, READ_WIDTH);
             #1 $finish;
           end
         case ({WRITE_P, READ_P})

             {"FALSE", "FALSE"} , {"TRUE", "TRUE"} :  ;

             {"FALSE", "TRUE"}: 
                begin 
                  $display("Port Width Mismatch on READ_WIDTH : The width READ_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  The parity bit(s) have not been written and hence cannot be read. ", READ_WIDTH);
                end
             {"TRUE", "FALSE"}: 
                begin 
                  $display("Port Width Mismatch on WRITE_WIDTH: The width WRITE_WIDTH on BRAM_SDP_MACRO instance %m is set to %d.  The parity bit(s) cannot be read ", WRITE_WIDTH);
	        end
          endcase
         
     end // end checks spartan6
    end // initial begin

   // Widths of Parity Bus
   localparam DIP_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (WRITE_WIDTH < 9) ? 0 : (WRITE_WIDTH == 9) ? 1 : (WRITE_WIDTH == 17) ? 1 : (WRITE_WIDTH == 18) ? 2 : (WRITE_WIDTH == 33) ? 1 : (WRITE_WIDTH == 34) ? 2 : (WRITE_WIDTH == 35) ? 3 : (WRITE_WIDTH == 36) ? 4 : (WRITE_WIDTH == 65) ? 1 : (WRITE_WIDTH == 66) ? 2 : (WRITE_WIDTH == 67) ? 3 : (WRITE_WIDTH == 68) ? 4 : (WRITE_WIDTH == 69) ? 5 : (WRITE_WIDTH == 70) ? 6 : (WRITE_WIDTH == 71) ? 7 : (WRITE_WIDTH == 72) ? 8 : 0 ) : 0;
  
   localparam DOP_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (READ_WIDTH < 9) ? 0 : (READ_WIDTH == 9) ? 1 : (READ_WIDTH == 17) ? 1 : (READ_WIDTH == 18) ? 2 : (READ_WIDTH == 33) ? 1 : (READ_WIDTH == 34) ? 2 : (READ_WIDTH == 35) ? 3 : (READ_WIDTH == 36) ? 4 : (READ_WIDTH == 65) ? 1 : (READ_WIDTH == 66) ? 2 : (READ_WIDTH == 67) ? 3 : (READ_WIDTH == 68) ? 4 : (READ_WIDTH == 69) ? 5 : (READ_WIDTH == 70) ? 6 : (READ_WIDTH == 71) ? 7 : (READ_WIDTH == 72) ? 8 : 0 ) : 0;

   // Widths of Data Bus
  localparam DI_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (WRITE_WIDTH == 1) ? 1 : (WRITE_WIDTH == 2) ? 2 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 4 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 8 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 16 : (BRAM_SIZE == "18Kb" && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? (WRITE_WIDTH-DIP_WIDTH) : (BRAM_SIZE == "36Kb" && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 32 : (BRAM_SIZE == "36Kb" && WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? (WRITE_WIDTH-DIP_WIDTH) : (WRITE_WIDTH-DIP_WIDTH) ): (WRITE_WIDTH-DIP_WIDTH);
  
  localparam DO_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (READ_WIDTH == 1) ? 1 : (READ_WIDTH == 2) ? 2 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 4 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 8 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 16 : (BRAM_SIZE == "18Kb" && READ_WIDTH > 18 && READ_WIDTH <= 36) ? (READ_WIDTH-DOP_WIDTH) : (BRAM_SIZE == "36Kb" && READ_WIDTH > 18 && READ_WIDTH <= 36) ? 32 : (BRAM_SIZE == "36Kb" && READ_WIDTH > 36 && READ_WIDTH <= 72) ? (READ_WIDTH-DOP_WIDTH) : (READ_WIDTH-DOP_WIDTH) ): (READ_WIDTH-DOP_WIDTH);

   // Widths of Address Bus
  localparam RDADDR_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (BRAM_SIZE == "9Kb") ? ( (READ_WIDTH == 1) ? 13 : (READ_WIDTH == 2) ? 12 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 11 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 10 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 9 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 8 : 13 ) : (BRAM_SIZE == "18Kb") ? ( (READ_WIDTH == 1) ? 14 : (READ_WIDTH == 2) ? 13 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 12 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 11 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 10 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 9 : 14 ) : (BRAM_SIZE == "36Kb") ? ( (READ_WIDTH == 1) ? 15 : (READ_WIDTH == 2) ? 14 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 13 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 12 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 11 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 10 : (READ_WIDTH > 36 && READ_WIDTH <= 72) ? 9 : 15 ) : 15) : 15;
  
  localparam WRADDR_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (BRAM_SIZE == "9Kb") ? ( (WRITE_WIDTH == 1) ? 13 : (WRITE_WIDTH == 2) ? 12 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 11 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 10 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 9 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 8 : 13 ) : (BRAM_SIZE == "18Kb") ? ( (WRITE_WIDTH == 1) ? 14 : (WRITE_WIDTH == 2) ? 13 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 12 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 11 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 10 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 9 : 14 ) : (BRAM_SIZE == "36Kb") ? ( (WRITE_WIDTH == 1) ? 15 : (WRITE_WIDTH == 2) ? 14 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 13 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 12 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 11 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 10 : (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? 9 : 15 ) : 15) : 15;
   // Widths of Write Enables
   localparam WE_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (WRITE_WIDTH <= 9) ? 1 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 2 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 4 : (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? 8 : (BRAM_SIZE == "18Kb") ? 4 : 8 ) : 8;
   
    localparam rd_width = (DEVICE == "VIRTEX5") ? ( (READ_WIDTH == 0) ? 0 : (READ_WIDTH == 1) ? 1 : (READ_WIDTH == 2) ? 2 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 4 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 9 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 18 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 36 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
  (DEVICE == "VIRTEX6" || DEVICE == "7SERIES") ? ( (READ_WIDTH == 0) ? 0 : (READ_WIDTH == 1) ? 1 : (READ_WIDTH == 2) ? 2 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 4 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 9 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 18 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 36 : (READ_WIDTH > 36 && READ_WIDTH <= 72) ? 72 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
  (DEVICE == "SPARTAN6") ? ( (READ_WIDTH == 0) ? 0 : (READ_WIDTH == 1) ? 1 : (READ_WIDTH == 2) ? 2 : (READ_WIDTH > 2 && READ_WIDTH <= 4) ? 4 : (READ_WIDTH > 4 && READ_WIDTH <= 9) ? 9 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 18 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 36 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
    36;

   localparam wr_width = (DEVICE == "VIRTEX5") ? ( (WRITE_WIDTH == 0) ? 0 : (WRITE_WIDTH == 1) ? 1 : (WRITE_WIDTH == 2) ? 2 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 4 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 9 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 18 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 36 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
    (DEVICE == "VIRTEX6" || DEVICE == "7SERIES") ? ( (WRITE_WIDTH == 0) ? 0 : (WRITE_WIDTH == 1) ? 1 : (WRITE_WIDTH == 2) ? 2 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 4 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 9 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 18 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 36 : (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? 72 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
    (DEVICE == "SPARTAN6") ? ( (WRITE_WIDTH == 0) ? 0 : (WRITE_WIDTH == 1) ? 1 : (WRITE_WIDTH == 2) ? 2 : (WRITE_WIDTH > 2 && WRITE_WIDTH <= 4) ? 4 : (WRITE_WIDTH > 4 && WRITE_WIDTH <= 9) ? 9 : (WRITE_WIDTH > 9 && WRITE_WIDTH <= 18) ? 18 : (WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 36 : (BRAM_SIZE == "18Kb") ? 18 : 36 ) :
   36;

localparam RD_BYTE_WIDTH = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (READ_WIDTH <= 9) ? 1 : (READ_WIDTH > 9 && READ_WIDTH <= 18) ? 2 : (READ_WIDTH > 18 && READ_WIDTH <= 36) ? 4 : (READ_WIDTH > 36 && READ_WIDTH <= 72) ? 8 : (BRAM_SIZE == "18Kb") ? 4 : 8 ) : 8;

localparam WR_WIDTHP = ((WRITE_WIDTH == 9) || (WRITE_WIDTH == 17) || (WRITE_WIDTH == 33) || (WRITE_WIDTH == 65)) ? 1 : ((WRITE_WIDTH == 18) || (WRITE_WIDTH == 34) || (WRITE_WIDTH == 66)) ? 2 : ((WRITE_WIDTH == 35) || (WRITE_WIDTH == 67)) ? 3 : ((WRITE_WIDTH == 36) || (WRITE_WIDTH == 68)) ? 4 : (WRITE_WIDTH == 69) ? 5 : (WRITE_WIDTH == 70) ? 6 : (WRITE_WIDTH == 71) ? 7 : (WRITE_WIDTH == 72) ? 8 : 8;

localparam RD_WIDTHP = ((READ_WIDTH == 9) || (READ_WIDTH == 17) || (READ_WIDTH == 33) || (READ_WIDTH == 65)) ? 1 : ((READ_WIDTH == 18) || (READ_WIDTH == 34) || (READ_WIDTH == 66)) ? 2 : ((READ_WIDTH == 35) || (READ_WIDTH == 67)) ? 3 : ((READ_WIDTH == 36) || (READ_WIDTH == 68)) ? 4 : (READ_WIDTH == 69) ? 5 : (READ_WIDTH == 70) ? 6 : (READ_WIDTH == 71) ? 7 : (READ_WIDTH == 72) ? 8 : 8;
   
   // Output Ports
   output [READ_WIDTH-1:0] DO;

   // Input Ports
   input [WRITE_WIDTH-1:0] DI;
   input RDCLK;
   input [RDADDR_WIDTH-1:0] RDADDR;
   input RDEN;
   input REGCE;
   input RST;
   input [WE_WIDTH-1:0] WE;
   input [WRADDR_WIDTH-1:0] WRADDR;
   input WRCLK;
   input WREN;

   // Mapping wire sizes _ for virtex5, read_width = write_width
   localparam greatest_width = (READ_WIDTH > WRITE_WIDTH) ? READ_WIDTH : WRITE_WIDTH;

   localparam MAX_ADDR_SIZE = (DEVICE == "VIRTEX5") ? ((BRAM_SIZE == "18Kb" && WRITE_WIDTH <= 18) ? 14 : (BRAM_SIZE == "18Kb" && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 9 : (BRAM_SIZE == "36Kb" && WRITE_WIDTH <= 36) ? 16 : (BRAM_SIZE == "36Kb" && WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? 9 : 16) :
  (DEVICE == "VIRTEX6" || DEVICE == "7SERIES") ? ( (BRAM_SIZE == "18Kb") ? 14 : 16 ) : 
  (DEVICE == "SPARTAN6") ? ( (BRAM_SIZE == "9Kb") ? 13 : 14 ) :
   16;
   localparam MAX_D_SIZE = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" ) ? ((BRAM_SIZE == "18Kb" && greatest_width <= 18) ? 16 : (BRAM_SIZE == "18Kb" && greatest_width > 18 && greatest_width <= 36) ? 32 : (BRAM_SIZE == "36Kb" && greatest_width <= 36) ? 32 : (BRAM_SIZE == "36Kb" && greatest_width > 36 && greatest_width <= 72) ? 64 : 64 ) :  
  (DEVICE == "SPARTAN6") ? ((BRAM_SIZE == "9Kb" && greatest_width <= 18) ? 16 : (BRAM_SIZE == "9Kb"  && greatest_width > 18 && greatest_width <= 36) ? 32 : 32 ) :
   32;
   localparam MAX_DP_SIZE = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" ) ? ( (BRAM_SIZE == "18Kb" && greatest_width <= 18) ? 2 : ( BRAM_SIZE == "18Kb" && greatest_width > 18 && greatest_width <= 36) ? 4 : (BRAM_SIZE == "36Kb" && greatest_width <= 36) ? 4 : ( BRAM_SIZE == "36Kb" && greatest_width > 36 && greatest_width <= 72) ? 8 : 8 ) : 
  (DEVICE == "SPARTAN6") ? ( (BRAM_SIZE == "9Kb" && greatest_width <= 18) ? 2 : (BRAM_SIZE == "9Kb"  && greatest_width > 18 && greatest_width <= 36) ? 4 : 4) :
   4;
   localparam MAX_WE_SIZE = (DEVICE == "VIRTEX5") ? ( (BRAM_SIZE == "18Kb" && WRITE_WIDTH <= 18) ? 2 : ( BRAM_SIZE == "18Kb" && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 4 : (BRAM_SIZE == "36Kb" && WRITE_WIDTH <= 36) ? 4 : ( BRAM_SIZE == "36Kb" && WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ? 8 : 8 ) :
   (DEVICE == "VIRTEX6" || DEVICE == "7SERIES") ? ( (BRAM_SIZE == "18Kb") ? 4 : 8 ) :
   (DEVICE == "SPARTAN6") ? ( (BRAM_SIZE == "9Kb"&& WRITE_WIDTH <= 18) ? 2 : (BRAM_SIZE == "9Kb"  && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) ? 4 : 4 ) :
    4;

   localparam fin_rd_width = (READ_WIDTH == 0) ? 1 : READ_WIDTH;
   localparam fin_wr_width = (WRITE_WIDTH == 0) ? 1 : WRITE_WIDTH;

   wire [MAX_ADDR_SIZE-1:0] RDADDR_PATTERN;
   wire [MAX_ADDR_SIZE-1:0] WRADDR_PATTERN;

   wire [MAX_ADDR_SIZE-1:0] RDADDR_PATTERN_SDP;
   wire [MAX_ADDR_SIZE-1:0] WRADDR_PATTERN_SDP;
   wire [MAX_D_SIZE-1:0] DI_PATTERN;
   wire [MAX_DP_SIZE-1:0] DIP_PATTERN;
   wire [MAX_D_SIZE-1:0] DO_PATTERN;
   wire [MAX_DP_SIZE-1:0] DOP_PATTERN;
   wire [MAX_WE_SIZE-1:0] WE_PATTERN;
   wire RSTRAM_PATTERN;
   wire RSTREG_PATTERN;

    // Pattern for WRADDR and RDADDR based on size of address  
   assign WRADDR_PATTERN  = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (BRAM_SIZE == "9Kb") ? ( (WRADDR_WIDTH == 13) ? WRADDR : (WRADDR_WIDTH == 12) ? {WRADDR, 1'b1} : (WRADDR_WIDTH == 11) ? {WRADDR, 2'b11} : (WRADDR_WIDTH == 10) ? {WRADDR, 3'b111} : (WRADDR_WIDTH == 9) ? {WRADDR, 4'b1111} : (WRADDR_WIDTH == 8) ? {WRADDR, 5'b11111} : WRADDR ) : (BRAM_SIZE == "18Kb") ? ( (WRADDR_WIDTH == 14) ? WRADDR : (WRADDR_WIDTH == 13) ? {WRADDR, 1'b1} : (WRADDR_WIDTH == 12) ? {WRADDR, 2'b11} : (WRADDR_WIDTH == 11) ? {WRADDR, 3'b111} : (WRADDR_WIDTH == 10) ? {WRADDR, 4'b1111} : (WRADDR_WIDTH == 9) ? {WRADDR, 5'b11111} : (WRADDR_WIDTH == 8) ? {WRADDR, 6'b111111} : WRADDR ) : (BRAM_SIZE == "36Kb") ? ( (WRADDR_WIDTH == 16) ? WRADDR : (WRADDR_WIDTH == 15) ? {1'b1, WRADDR} : (WRADDR_WIDTH == 14) ? {1'b1, WRADDR, 1'b1} : (WRADDR_WIDTH == 13) ? {1'b1, WRADDR, 2'b11} : (WRADDR_WIDTH == 12) ? {1'b1, WRADDR, 3'b111} : (WRADDR_WIDTH == 11) ? {1'b1, WRADDR, 4'b1111} : (WRADDR_WIDTH == 10) ? {1'b1, WRADDR, 5'b11111} : (WRADDR_WIDTH == 9) ? {1'b1, WRADDR, 6'b111111}  : WRADDR ) : WRADDR ) : WRADDR;

   assign RDADDR_PATTERN  = (DEVICE == "VIRTEX5" || DEVICE == "VIRTEX6" || DEVICE == "7SERIES" || DEVICE == "SPARTAN6" ) ? ( (BRAM_SIZE == "9Kb") ? ( (RDADDR_WIDTH == 13) ? RDADDR : (RDADDR_WIDTH == 12) ? {RDADDR, 1'b1} : (RDADDR_WIDTH == 11) ? {RDADDR, 2'b11} : (RDADDR_WIDTH == 10) ? {RDADDR, 3'b111} : (RDADDR_WIDTH == 9) ? {RDADDR, 4'b1111} : (RDADDR_WIDTH == 8) ? {RDADDR, 5'b11111} : RDADDR ) : (BRAM_SIZE == "18Kb") ? ( (RDADDR_WIDTH == 14) ? RDADDR : (RDADDR_WIDTH == 13) ? {RDADDR, 1'b1} : (RDADDR_WIDTH == 12) ? {RDADDR, 2'b11} : (RDADDR_WIDTH == 11) ? {RDADDR, 3'b111} : (RDADDR_WIDTH == 10) ? {RDADDR, 4'b1111} : (RDADDR_WIDTH == 9) ? {RDADDR, 5'b11111} : (RDADDR_WIDTH == 8) ? {RDADDR, 6'b11111} : RDADDR ) : (BRAM_SIZE == "36Kb") ? ( (RDADDR_WIDTH == 16) ? RDADDR : (RDADDR_WIDTH == 15) ? {1'b1, RDADDR} : (RDADDR_WIDTH == 14) ? {1'b1, RDADDR, 1'b1} : (RDADDR_WIDTH == 13) ? {1'b1, RDADDR, 2'b11} : (RDADDR_WIDTH == 12) ? {1'b1, RDADDR, 3'b111} : (RDADDR_WIDTH == 11) ? {1'b1, RDADDR, 4'b1111} : (RDADDR_WIDTH == 10) ? {1'b1, RDADDR, 5'b11111} : (RDADDR_WIDTH == 9) ? {1'b1, RDADDR, 6'b111111}  : RDADDR ) : RDADDR ) : RDADDR;
    
   localparam INIT_SRVAL_WIDTH_SIZE = (BRAM_SIZE == "36Kb") ? ((READ_WIDTH > 36 || WRITE_WIDTH > 36) ? 72 : 36) : 
				      (BRAM_SIZE == "18Kb") ? ((DEVICE == "SPARTAN6" || (READ_WIDTH > 18 || WRITE_WIDTH > 18)) ? 36 : 18) : 
				      (BRAM_SIZE == "9Kb") ? ((WRITE_WIDTH > 18) ? 36 : 18) : 36;
   
   localparam init_tmp = (READ_P == "TRUE" && WRITE_P == "TRUE") ? 
			 ((READ_WIDTH == 9) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {9'b0,INIT[8],INIT[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {27'b0,INIT[8],INIT[7:0]} : {63'b0,INIT[8],INIT[7:0]}) :
			  (READ_WIDTH == 17) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {1'b0,INIT[8],INIT[16:9],INIT[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {19'b0,INIT[8],INIT[16:9],INIT[7:0]} : {55'b0,INIT[8],INIT[16:9],INIT[7:0]}) :
			  (READ_WIDTH == 18) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {INIT[17],INIT[8],INIT[16:9],INIT[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {18'b0,INIT[17],INIT[8],INIT[16:9],INIT[7:0]} : {54'b0,INIT[17],INIT[8],INIT[16:9],INIT[7:0]}) :
			  (READ_WIDTH == 33) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {3'b0,INIT[8],INIT[32:9],INIT[7:0]} : {39'b0,INIT[8],INIT[32:9],INIT[7:0]}) :
			  (READ_WIDTH == 34) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {2'b0,INIT[17],INIT[8],INIT[33:18],INIT[16:9],INIT[7:0]} : {38'b0,INIT[17],INIT[8],INIT[33:18],INIT[16:9],INIT[7:0]}) :
			  (READ_WIDTH == 35) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {1'b0,INIT[26],INIT[17],INIT[8],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} : {37'b0,INIT[26],INIT[17],INIT[8],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]}) :
 			  (READ_WIDTH == 36) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {INIT[35],INIT[26],INIT[17],INIT[8],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} : {36'b0,INIT[35],INIT[26],INIT[17],INIT[8],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]}) :
                          (READ_WIDTH == 65) ? {7'b0,INIT[8],INIT[64:9],INIT[7:0]} :
			  (READ_WIDTH == 66) ? {6'b0,INIT[17],INIT[8],INIT[65:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 67) ? {5'b0,INIT[26],INIT[17],INIT[8],INIT[66:27],INIT[25:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 68) ? {4'b0,INIT[35],INIT[26],INIT[17],INIT[8],INIT[67:36],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 69) ? {3'b0,INIT[44],INIT[35],INIT[26],INIT[17],INIT[8],INIT[68:45],INIT[43:36],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 70) ? {2'b0,INIT[53],INIT[44],INIT[35],INIT[26],INIT[17],INIT[8],INIT[69:54],INIT[52:45],INIT[43:36],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 71) ? {1'b0,INIT[62],INIT[53],INIT[44],INIT[35],INIT[26],INIT[17],INIT[8],INIT[70:63],INIT[61:54],INIT[52:45],INIT[43:36],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} :
			  (READ_WIDTH == 72) ? {INIT[71],INIT[62],INIT[53],INIT[44],INIT[35],INIT[26],INIT[17],INIT[8],INIT[70:63],INIT[61:54],INIT[52:45],INIT[43:36],INIT[34:27],INIT[25:18],INIT[16:9],INIT[7:0]} : INIT) : INIT;		  


   localparam srval_tmp = (READ_P == "TRUE" && WRITE_P == "TRUE") ? 
			 ((READ_WIDTH == 9) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {9'b0,SRVAL[8],SRVAL[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {27'b0,SRVAL[8],SRVAL[7:0]} : {63'b0,SRVAL[8],SRVAL[7:0]}) :
			  (READ_WIDTH == 17) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {1'b0,SRVAL[8],SRVAL[16:9],SRVAL[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {19'b0,SRVAL[8],SRVAL[16:9],SRVAL[7:0]} : {55'b0,SRVAL[8],SRVAL[16:9],SRVAL[7:0]}) :
			  (READ_WIDTH == 18) ? ((INIT_SRVAL_WIDTH_SIZE == 18) ? {SRVAL[17],SRVAL[8],SRVAL[16:9],SRVAL[7:0]} : (INIT_SRVAL_WIDTH_SIZE == 36) ? {18'b0,SRVAL[17],SRVAL[8],SRVAL[16:9],SRVAL[7:0]} : {54'b0,SRVAL[17],SRVAL[8],SRVAL[16:9],SRVAL[7:0]}) :
			  (READ_WIDTH == 33) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {3'b0,SRVAL[8],SRVAL[32:9],SRVAL[7:0]} : {39'b0,SRVAL[8],SRVAL[32:9],SRVAL[7:0]}) :
			  (READ_WIDTH == 34) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {2'b0,SRVAL[17],SRVAL[8],SRVAL[33:18],SRVAL[16:9],SRVAL[7:0]} : {38'b0,SRVAL[17],SRVAL[8],SRVAL[33:18],SRVAL[16:9],SRVAL[7:0]}) :
			  (READ_WIDTH == 35) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {1'b0,SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} : {37'b0,SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]}) :
 			  (READ_WIDTH == 36) ? ((INIT_SRVAL_WIDTH_SIZE == 36) ? {SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} : {36'b0,SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]}) :
                          (READ_WIDTH == 65) ? {7'b0,SRVAL[8],SRVAL[64:9],SRVAL[7:0]} :
			  (READ_WIDTH == 66) ? {6'b0,SRVAL[17],SRVAL[8],SRVAL[65:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 67) ? {5'b0,SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[66:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 68) ? {4'b0,SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[67:36],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 69) ? {3'b0,SRVAL[44],SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[68:45],SRVAL[43:36],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 70) ? {2'b0,SRVAL[53],SRVAL[44],SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[69:54],SRVAL[52:45],SRVAL[43:36],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 71) ? {1'b0,SRVAL[62],SRVAL[53],SRVAL[44],SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[70:63],SRVAL[61:54],SRVAL[52:45],SRVAL[43:36],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} :
			  (READ_WIDTH == 72) ? {SRVAL[71],SRVAL[62],SRVAL[53],SRVAL[44],SRVAL[35],SRVAL[26],SRVAL[17],SRVAL[8],SRVAL[70:63],SRVAL[61:54],SRVAL[52:45],SRVAL[43:36],SRVAL[34:27],SRVAL[25:18],SRVAL[16:9],SRVAL[7:0]} : SRVAL) : SRVAL;
   
   
   genvar i, i1, j, j1, j2;
   wire [DIP_WIDTH-1:0] DIP_tmp = 'b0;
   
  // Pattern for DATA bus
    generate
      case(DEVICE)
        "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6" : 
	   if ( (BRAM_SIZE == "9Kb" && READ_WIDTH <= 36) || (BRAM_SIZE == "18Kb" && READ_WIDTH <= 36) || (BRAM_SIZE == "36Kb" && READ_WIDTH <= 72))
             begin : di1
		if ((READ_P == "TRUE" && WRITE_P == "TRUE") && ( (BRAM_SIZE == "9Kb" && WRITE_WIDTH == 36) || (BRAM_SIZE == "18Kb" && WRITE_WIDTH == 36) || (BRAM_SIZE == "36Kb" && WRITE_WIDTH == 72)))
                begin : di1

		   if (WRITE_WIDTH >= 71 || WRITE_WIDTH == 35 || WRITE_WIDTH == 36 || WRITE_WIDTH <= 32) begin : di221
		      for (i = 0; i < WE_WIDTH; i = i + 1) begin : di_byte1
			 assign DI_PATTERN[(i*8) +: 8] = DI[((i*8)+i) +: 8];
		      end
		   end
		   
		   if (WRITE_WIDTH == 33) begin : di222
		      assign DI_PATTERN = {DI[32:9], DI[7:0]};
		   end
		   
		   if (WRITE_WIDTH == 34) begin : di223
		      assign DI_PATTERN = {DI[33:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 65) begin : di224
		      assign DI_PATTERN = {DI[64:9], DI[7:0]};
		   end
		   
		   if (WRITE_WIDTH == 66) begin : di225
		      assign DI_PATTERN = {DI[65:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 67) begin : di226
		      assign DI_PATTERN = {DI[66:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end
		   
		   if (WRITE_WIDTH == 68) begin : di227
		      assign DI_PATTERN = {DI[67:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 69) begin : di228
		      assign DI_PATTERN = {DI[68:45], DI[43:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 70) begin : di229
		      assign DI_PATTERN = {DI[69:54], DI[52:45], DI[43:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   for (j = 1; j <= WR_WIDTHP; j = j + 1) begin : dip_byte1
		     assign DIP_PATTERN[j-1] = DI[((j*8)+j-1)];
		   end
                end
	        else if ((READ_P == "TRUE" && WRITE_P == "TRUE") && ( (BRAM_SIZE == "9Kb" && WRITE_WIDTH < 36) || (BRAM_SIZE == "18Kb" && WRITE_WIDTH < 36) || (BRAM_SIZE == "36Kb" && WRITE_WIDTH < 72)))
		begin : di2 

		   if (WRITE_WIDTH >= 71 || WRITE_WIDTH == 35 || WRITE_WIDTH == 36 || WRITE_WIDTH <= 32) begin : di221
		      for (i = 0; i < WE_WIDTH; i = i + 1) begin : di_byte2
			 assign DI_PATTERN[(i*8) +: 8] = DI[((i*8)+i) +: 8];
		      end
		   end
		   
		   if (WRITE_WIDTH == 33) begin : di222
		      assign DI_PATTERN = {DI[32:9], DI[7:0]};
		   end
	       
		   if (WRITE_WIDTH == 34) begin : di223
		      assign DI_PATTERN = {DI[33:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 65) begin : di224
		      assign DI_PATTERN = {DI[64:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 66) begin : di225
		      assign DI_PATTERN = {DI[65:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 67) begin : di226
		      assign DI_PATTERN = {DI[66:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 68) begin : di227
		      assign DI_PATTERN = {DI[67:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 69) begin : di228
		      assign DI_PATTERN = {DI[68:45], DI[43:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end

		   if (WRITE_WIDTH == 70) begin : di229
		      assign DI_PATTERN = {DI[69:54], DI[52:45], DI[43:36], DI[34:27], DI[25:18],  DI[16:9], DI[7:0]};
		   end


		   for (j = 1; j <= WR_WIDTHP; j = j + 1) begin : dip_byte2
		      assign DIP_PATTERN[j-1] = DI[((j*8)+j-1)];
		   end
		   
		   for (j2 = DIP_WIDTH; j2 < MAX_DP_SIZE; j2 = j2 + 1) begin : dip_byte2_0
		      assign DIP_PATTERN[j2] = 1'b0;
		   end
		   
		end
                else if ( (READ_P == "FALSE" && WRITE_P == "FALSE") && ( (BRAM_SIZE == "9Kb" && WRITE_WIDTH == 32) || (BRAM_SIZE == "18Kb" && WRITE_WIDTH == 32) || (BRAM_SIZE == "36Kb" && WRITE_WIDTH == 64)))
                begin : di3
                   assign DI_PATTERN = DI;
                   assign DIP_PATTERN = 0;
                end
	        else if ( (READ_P == "FALSE" && WRITE_P == "FALSE") && ((READ_WIDTH == WRITE_WIDTH) || (READ_WIDTH/WRITE_WIDTH == 2) || (valid_width == "TRUE")) )	
		begin : di4
                   assign DI_PATTERN = {{((MAX_D_SIZE)-fin_wr_width){1'b0}}, DI};
		   assign DIP_PATTERN = 0;
                end
                else if ( (READ_WIDTH == 1 && WRITE_WIDTH == 2) || (READ_WIDTH == 2 && WRITE_WIDTH == 4) || (READ_WIDTH == 4 && WRITE_WIDTH == 8) || (READ_WIDTH == 8 && WRITE_WIDTH == 16)|| (READ_WIDTH == 16 && WRITE_WIDTH == 32)|| (READ_WIDTH == 32 && WRITE_WIDTH == 64 ) )
		begin : dird
		   assign DI_PATTERN = {{((MAX_D_SIZE)-fin_wr_width){1'b0}}, DI};
		end
		else if ( (READ_P == "FALSE" && WRITE_P == "FALSE") && (WRITE_WIDTH/READ_WIDTH == 2))
		begin
		  if (READ_WIDTH == 3)
	            begin : dird3
		       assign DI_PATTERN = { {{(4-READ_WIDTH)}{1'b0}}, DI[((2*READ_WIDTH)-1):READ_WIDTH], {{(4-READ_WIDTH)}{1'b0}}, DI[(READ_WIDTH-1):0]};
		    end
		    else if (READ_WIDTH > 4 && READ_WIDTH < 8)
		    begin : dird567
		       assign DI_PATTERN = { {{(8-READ_WIDTH)}{1'b0}}, DI[((2*READ_WIDTH)-1):READ_WIDTH], {{(8-READ_WIDTH)}{1'b0}}, DI[(READ_WIDTH-1):0]};
		    end
		    else if (READ_WIDTH > 8 && READ_WIDTH < 16)
		    begin : dird915
		       assign DI_PATTERN = { {{(16-READ_WIDTH)}{1'b0}}, DI[((2*READ_WIDTH)-1):READ_WIDTH], {{(16-READ_WIDTH)}{1'b0}} ,DI[(READ_WIDTH-1):0]};
		    end   
		    else if (READ_WIDTH > 16 && READ_WIDTH < 32)
		    begin : dird1632
		       assign DI_PATTERN = { {{(32-READ_WIDTH)}{1'b0}}, DI[((2*READ_WIDTH)-1):READ_WIDTH], {{(32-READ_WIDTH)}{1'b0}}, DI[(READ_WIDTH-1):0]};
		    end     
		    else
		    begin
		       assign DI_PATTERN = {{((MAX_D_SIZE)-fin_wr_width){1'b0}}, DI};
		    end
		 end   
           end
      endcase
   endgenerate
   generate 
      case(DEVICE)
        "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6" : 
           if ( (BRAM_SIZE == "9Kb" && READ_WIDTH <= 36) || (BRAM_SIZE == "18Kb" && READ_WIDTH <= 36) || (BRAM_SIZE == "36Kb" && READ_WIDTH <= 72))
	     begin : do1
	        if ((READ_P == "TRUE") && (WRITE_P == "TRUE"))
		begin : do11

		   if (READ_WIDTH >= 71 || READ_WIDTH == 35 || READ_WIDTH == 36 || READ_WIDTH <= 32) begin : do_byte11
		      for (i1 = 0; i1 < RD_BYTE_WIDTH; i1 = i1 + 1) begin : do_byte1
			 assign DO[((i1*8)+i1) +: 8] = DO_PATTERN[(i1*8) +: 8];
		      end
		   end

		   if (READ_WIDTH == 33) begin : do_byte12
		      assign DO[32:9] = DO_PATTERN[31:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end
		   
		   if (READ_WIDTH == 34) begin : do_byte13
		      assign DO[33:18] = DO_PATTERN[31:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end
		   
		   if (READ_WIDTH == 65) begin : do_byte14
		      assign DO[64:9] = DO_PATTERN[63:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   if (READ_WIDTH == 66) begin : do_byte15
		      assign DO[65:18] = DO_PATTERN[63:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   if (READ_WIDTH == 67) begin : do_byte16
		      assign DO[66:27] = DO_PATTERN[63:24];
		      assign DO[25:18] = DO_PATTERN[23:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   if (READ_WIDTH == 68) begin : do_byte17
		      assign DO[67:36] = DO_PATTERN[63:32];
		      assign DO[34:27] = DO_PATTERN[31:24];
		      assign DO[25:18] = DO_PATTERN[23:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   if (READ_WIDTH == 69) begin : do_byte18
		      assign DO[68:45] = DO_PATTERN[63:40];
		      assign DO[43:36] = DO_PATTERN[39:32];
		      assign DO[34:27] = DO_PATTERN[31:24];
		      assign DO[25:18] = DO_PATTERN[23:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   if (READ_WIDTH == 70) begin : do_byte19
		      assign DO[69:54] = DO_PATTERN[63:48];
		      assign DO[52:45] = DO_PATTERN[47:40];
		      assign DO[43:36] = DO_PATTERN[39:32];
		      assign DO[34:27] = DO_PATTERN[31:24];
		      assign DO[25:18] = DO_PATTERN[23:16];
		      assign DO[16:9] = DO_PATTERN[15:8];
		      assign DO[7:0] = DO_PATTERN[7:0];
		   end

		   
		   for (j1 = 1; j1 <= RD_WIDTHP; j1 = j1 + 1) begin : dop_byte1
		     assign DO[((j1*8)+j1-1)] = DOP_PATTERN[j1-1];
		   end
		   
		   
                end
		else if ( (READ_P == "FALSE" && WRITE_P == "FALSE") && ((READ_WIDTH == WRITE_WIDTH) || (WRITE_WIDTH/READ_WIDTH == 2) || (valid_width == "TRUE")) )
		begin : do2
                  assign DO = DO_PATTERN[fin_rd_width-1:0];
		end
		else if ( (READ_WIDTH == 2 && WRITE_WIDTH == 1) || (READ_WIDTH == 4 && WRITE_WIDTH == 2) || (READ_WIDTH == 8 && WRITE_WIDTH == 4) || (READ_WIDTH == 16 && WRITE_WIDTH == 8)|| (READ_WIDTH == 32 && WRITE_WIDTH == 16)|| (READ_WIDTH == 64 && WRITE_WIDTH == 32 ) )
		begin
		     assign DO = DO_PATTERN[fin_rd_width-1:0];
		end
		else if ( (READ_P == "FALSE" && WRITE_P == "FALSE") && (READ_WIDTH/WRITE_WIDTH == 2))
		begin
		    if (WRITE_WIDTH == 3)
	            begin : dowr3
		          assign DO = {DO_PATTERN[(4+(WRITE_WIDTH-1)):4], DO_PATTERN[(WRITE_WIDTH-1):0]};
		    end
		    else if (WRITE_WIDTH > 4 && WRITE_WIDTH < 8)
		    begin : dowr567
		        assign DO = {DO_PATTERN[(8+(WRITE_WIDTH-1)):8], DO_PATTERN[(WRITE_WIDTH-1):0]};
		    end
		    else if (WRITE_WIDTH > 8 && WRITE_WIDTH < 16)
		    begin : dowr915
		        assign DO = {DO_PATTERN[(16+(WRITE_WIDTH-1)):16], DO_PATTERN[(WRITE_WIDTH-1):0]};
		    end   
		    else if (WRITE_WIDTH > 16 && WRITE_WIDTH < 32)
		    begin : dowr1632
		        assign DO = {DO_PATTERN[(32+(WRITE_WIDTH-1)):32], DO_PATTERN[(WRITE_WIDTH-1):0]};
		    end     
		    else
		    begin
		    assign DO = DO_PATTERN[fin_rd_width-1:0];
		    end
		 end   
           end
      endcase
   endgenerate

   assign WE_PATTERN =  (BRAM_SIZE == "9Kb") ? ( (WE_WIDTH == 1) ? {2{WE}} : (WE_WIDTH == 2) ? WE : WE) : (BRAM_SIZE == "18Kb") ? ( (WE_WIDTH == 1) ? {4{WE}} : (WE_WIDTH == 2) ? {2{WE}} : (WE_WIDTH == 4) ? WE : WE) : (BRAM_SIZE == "36Kb") ? ( (WE_WIDTH == 1) ? {8{WE}} : (WE_WIDTH == 2) ? {4{WE}} : (WE_WIDTH == 4) ? {2{WE}} :(WE_WIDTH == 8) ? WE : WE) : WE;

   assign RSTREG_PATTERN = (DO_REG == 1'b1) ? RST : 1'b0; 
   assign RSTRAM_PATTERN = RST;
 
   localparam sim_device_pm = (DEVICE == "VIRTEX6") ? "VIRTEX6" : "7SERIES";
 
    generate 
      case(DEVICE)
        "VIRTEX5" : 
           begin
             if (BRAM_SIZE == "18Kb" && WRITE_WIDTH <= 18) begin : bram18_dp
              RAMB18 # ( 
                .DOA_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A (init_tmp),
                .INIT_B (init_tmp),
                .INIT_FILE(INIT_FILE),
                .READ_WIDTH_A (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_MODE (SIM_MODE),
                .SRVAL_A (srval_tmp),
                .WRITE_MODE_B ("READ_FIRST"),
                .WRITE_WIDTH_B (wr_width)
                )  bram18_tdp (
                .DOA (DO_PATTERN), 
                .DOB (), 
                .DOPA (DOP_PATTERN), 
                .DOPB (),
                .ADDRA(RDADDR_PATTERN), 
                .ADDRB(WRADDR_PATTERN), 
                .CLKA (RDCLK), 
                .CLKB (WRCLK), 
                .DIA (16'b0), 
                .DIB (DI_PATTERN), 
                .DIPA (2'b0), 
                .DIPB (DIP_PATTERN), 
                .ENA (RDEN), 
                .ENB (WREN), 
                .REGCEA (REGCE), 
                .REGCEB (1'b0), 
                .SSRA (RST), 
                .SSRB (1'b0), 
                .WEA (2'b0), 
                .WEB (WE_PATTERN)
                );
              end
             else if (BRAM_SIZE == "18Kb" && (WRITE_WIDTH > 18 && WRITE_WIDTH <=36)) begin : bram18_sdp
   
             RAMB18SDP # (
               .DO_REG (DO_REG), 
               .INIT (init_tmp),
               .INITP_00 (INITP_00),
               .INITP_01 (INITP_01),
               .INITP_02 (INITP_02), 
               .INITP_03 (INITP_03),
               .INITP_04 (INITP_04),
               .INITP_05 (INITP_05),
               .INITP_06 (INITP_06),
               .INITP_07 (INITP_07),
               .INIT_00 (INIT_00), 
               .INIT_01 (INIT_01),
               .INIT_02 (INIT_02),
               .INIT_03 (INIT_03),
               .INIT_04 (INIT_04),
               .INIT_05 (INIT_05),
               .INIT_06 (INIT_06),
               .INIT_07 (INIT_07),
               .INIT_08 (INIT_08),
               .INIT_09 (INIT_09),
               .INIT_0A (INIT_0A),
               .INIT_0B (INIT_0B),
               .INIT_0C (INIT_0C),
               .INIT_0D (INIT_0D),
               .INIT_0E (INIT_0E),
               .INIT_0F (INIT_0F),
               .INIT_10 (INIT_10),
               .INIT_11 (INIT_11),
               .INIT_12 (INIT_12),
               .INIT_13 (INIT_13),
               .INIT_14 (INIT_14),
               .INIT_15 (INIT_15),
               .INIT_16 (INIT_16),
               .INIT_17 (INIT_17),
               .INIT_18 (INIT_18),
               .INIT_19 (INIT_19),
               .INIT_1A (INIT_1A),
               .INIT_1B (INIT_1B),
               .INIT_1C (INIT_1C),
               .INIT_1D (INIT_1D),
               .INIT_1E (INIT_1E),
               .INIT_1F (INIT_1F),
               .INIT_20 (INIT_20),
               .INIT_21 (INIT_21),
               .INIT_22 (INIT_22),
               .INIT_23 (INIT_23),
               .INIT_24 (INIT_24),
               .INIT_25 (INIT_25),
               .INIT_26 (INIT_26),
               .INIT_27 (INIT_27),
               .INIT_28 (INIT_28),
               .INIT_29 (INIT_29),
               .INIT_2A (INIT_2A),
               .INIT_2B (INIT_2B),
               .INIT_2C (INIT_2C),
               .INIT_2D (INIT_2D),
               .INIT_2E (INIT_2E),
               .INIT_2F (INIT_2F),
               .INIT_30 (INIT_30),
               .INIT_31 (INIT_31),
               .INIT_32 (INIT_32),
               .INIT_33 (INIT_33),
               .INIT_34 (INIT_34),
               .INIT_35 (INIT_35),
               .INIT_36 (INIT_36),
               .INIT_37 (INIT_37),
               .INIT_38 (INIT_38),
               .INIT_39 (INIT_39),
               .INIT_3A (INIT_3A),
               .INIT_3B (INIT_3B),
               .INIT_3C (INIT_3C),
               .INIT_3D (INIT_3D),
               .INIT_3E (INIT_3E),
               .INIT_3F (INIT_3F),
               .INIT_FILE (INIT_FILE),
               .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
               .SIM_MODE (SIM_MODE),
               .SRVAL(srval_tmp) 
               ) bram18_sdp (
               .DO (DO_PATTERN), 
               .DOP (DOP_PATTERN), 
               .DI (DI_PATTERN), 
               .DIP (DIP_PATTERN), 
               .RDADDR (RDADDR), 
               .RDCLK (RDCLK), 
               .RDEN (RDEN), 
               .REGCE (REGCE), 
               .SSR (RST),  
               .WE (WE_PATTERN), 
               .WRADDR (WRADDR), 
               .WRCLK (WRCLK), 
               .WREN (WREN)
               );
            end 
          else if (BRAM_SIZE == "36Kb" && WRITE_WIDTH <= 36) begin : bram36_dp
   
          RAMB36 # ( 
              .DOA_REG (DO_REG),
              .INITP_00 (INITP_00),
              .INITP_01 (INITP_01),
              .INITP_02 (INITP_02), 
              .INITP_03 (INITP_03),
              .INITP_04 (INITP_04),
              .INITP_05 (INITP_05),
              .INITP_06 (INITP_06),
              .INITP_07 (INITP_07),
              .INIT_00 (INIT_00), 
              .INIT_01 (INIT_01),
              .INIT_02 (INIT_02),
              .INIT_03 (INIT_03),
              .INIT_04 (INIT_04),
              .INIT_05 (INIT_05),
              .INIT_06 (INIT_06),
              .INIT_07 (INIT_07),
              .INIT_08 (INIT_08),
              .INIT_09 (INIT_09),
              .INIT_0A (INIT_0A),
              .INIT_0B (INIT_0B),
              .INIT_0C (INIT_0C),
              .INIT_0D (INIT_0D),
              .INIT_0E (INIT_0E),
              .INIT_0F (INIT_0F),
              .INIT_10 (INIT_10),
              .INIT_11 (INIT_11),
              .INIT_12 (INIT_12),
              .INIT_13 (INIT_13),
              .INIT_14 (INIT_14),
              .INIT_15 (INIT_15),
              .INIT_16 (INIT_16),
              .INIT_17 (INIT_17),
              .INIT_18 (INIT_18),
              .INIT_19 (INIT_19),
              .INIT_1A (INIT_1A),
              .INIT_1B (INIT_1B),
              .INIT_1C (INIT_1C),
              .INIT_1D (INIT_1D),
              .INIT_1E (INIT_1E),
              .INIT_1F (INIT_1F),
              .INIT_20 (INIT_20),
              .INIT_21 (INIT_21),
              .INIT_22 (INIT_22),
              .INIT_23 (INIT_23),
              .INIT_24 (INIT_24),
              .INIT_25 (INIT_25),
              .INIT_26 (INIT_26),
              .INIT_27 (INIT_27),
              .INIT_28 (INIT_28),
              .INIT_29 (INIT_29),
              .INIT_2A (INIT_2A),
              .INIT_2B (INIT_2B),
              .INIT_2C (INIT_2C),
              .INIT_2D (INIT_2D),
              .INIT_2E (INIT_2E),
              .INIT_2F (INIT_2F),
              .INIT_30 (INIT_30),
              .INIT_31 (INIT_31),
              .INIT_32 (INIT_32),
              .INIT_33 (INIT_33),
              .INIT_34 (INIT_34),
              .INIT_35 (INIT_35),
              .INIT_36 (INIT_36),
              .INIT_37 (INIT_37),
              .INIT_38 (INIT_38),
              .INIT_39 (INIT_39),
              .INIT_3A (INIT_3A),
              .INIT_3B (INIT_3B),
              .INIT_3C (INIT_3C),
              .INIT_3D (INIT_3D),
              .INIT_3E (INIT_3E),
              .INIT_3F (INIT_3F),
              .INIT_40 (INIT_40), 
              .INIT_41 (INIT_41),
              .INIT_42 (INIT_42),
              .INIT_43 (INIT_43),
              .INIT_44 (INIT_44),
              .INIT_45 (INIT_45),
              .INIT_46 (INIT_46),
              .INIT_47 (INIT_47),
              .INIT_48 (INIT_48),
              .INIT_49 (INIT_49),
              .INIT_4A (INIT_4A),
              .INIT_4B (INIT_4B),
              .INIT_4C (INIT_4C),
              .INIT_4D (INIT_4D),
              .INIT_4E (INIT_4E),
              .INIT_4F (INIT_4F),
              .INIT_50 (INIT_50),
              .INIT_51 (INIT_51),
              .INIT_52 (INIT_52),
              .INIT_53 (INIT_53),
              .INIT_54 (INIT_54),
              .INIT_55 (INIT_55),
              .INIT_56 (INIT_56),
              .INIT_57 (INIT_57),
              .INIT_58 (INIT_58),
              .INIT_59 (INIT_59),
              .INIT_5A (INIT_5A),
              .INIT_5B (INIT_5B),
              .INIT_5C (INIT_5C),
              .INIT_5D (INIT_5D),
              .INIT_5E (INIT_5E),
              .INIT_5F (INIT_5F),
              .INIT_60 (INIT_60),
              .INIT_61 (INIT_61),
              .INIT_62 (INIT_62),
              .INIT_63 (INIT_63),
              .INIT_64 (INIT_64),
              .INIT_65 (INIT_65),
              .INIT_66 (INIT_66),
              .INIT_67 (INIT_67),
              .INIT_68 (INIT_68),
              .INIT_69 (INIT_69),
              .INIT_6A (INIT_6A),
              .INIT_6B (INIT_6B),
              .INIT_6C (INIT_6C),
              .INIT_6D (INIT_6D),
              .INIT_6E (INIT_6E),
              .INIT_6F (INIT_6F),
              .INIT_70 (INIT_70),
              .INIT_71 (INIT_71),
              .INIT_72 (INIT_72),
              .INIT_73 (INIT_73),
              .INIT_74 (INIT_74),
              .INIT_75 (INIT_75),
              .INIT_76 (INIT_76),
              .INIT_77 (INIT_77),
              .INIT_78 (INIT_78),
              .INIT_79 (INIT_79),
              .INIT_7A (INIT_7A),
              .INIT_7B (INIT_7B),
              .INIT_7C (INIT_7C),
              .INIT_7D (INIT_7D),
              .INIT_7E (INIT_7E),
              .INIT_7F (INIT_7F),
              .INIT_A (init_tmp),
              .INIT_FILE (INIT_FILE),
              .READ_WIDTH_A (rd_width),
              .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
              .SIM_MODE (SIM_MODE),
              .SRVAL_A (srval_tmp),
              .WRITE_MODE_B ("READ_FIRST"),
              .WRITE_WIDTH_B (wr_width)
              )  bram36_tdp (
              .CASCADEOUTLATA (),
              .CASCADEOUTLATB (),
              .CASCADEOUTREGA (),
              .CASCADEOUTREGB (),
              .DOA (DO_PATTERN), 
              .DOB (), 
              .DOPA (DOP_PATTERN), 
              .DOPB (),
              .ADDRA (RDADDR_PATTERN), 
              .ADDRB (WRADDR_PATTERN),
              .CASCADEINLATA (1'b0),
              .CASCADEINLATB (1'b0),
              .CASCADEINREGA (1'b0),
              .CASCADEINREGB (1'b0), 
              .CLKA (RDCLK), 
              .CLKB (WRCLK), 
              .DIA (32'b0), 
              .DIB (DI_PATTERN), 
              .DIPA (4'b0), 
              .DIPB (DIP_PATTERN), 
              .ENA (RDEN), 
              .ENB (WREN), 
              .REGCEA (REGCE), 
              .REGCEB (1'b0), 
              .SSRA (RST), 
              .SSRB (1'b0), 
              .WEA (4'b0), 
              .WEB (WE_PATTERN)
              );
            end

            else if (BRAM_SIZE == "36Kb" && (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72)) begin : bram36_sdp
   
            RAMB36SDP # (
               .DO_REG (DO_REG), 
               .INIT (init_tmp),
               .INITP_00 (INITP_00),
               .INITP_01 (INITP_01),
               .INITP_02 (INITP_02), 
               .INITP_03 (INITP_03),
               .INITP_04 (INITP_04),
               .INITP_05 (INITP_05),
               .INITP_06 (INITP_06),
               .INITP_07 (INITP_07),
               .INIT_00 (INIT_00), 
               .INIT_01 (INIT_01),
               .INIT_02 (INIT_02),
               .INIT_03 (INIT_03),
               .INIT_04 (INIT_04),
               .INIT_05 (INIT_05),
               .INIT_06 (INIT_06),
               .INIT_07 (INIT_07),
               .INIT_08 (INIT_08),
               .INIT_09 (INIT_09),
               .INIT_0A (INIT_0A),
               .INIT_0B (INIT_0B),
               .INIT_0C (INIT_0C),
               .INIT_0D (INIT_0D),
               .INIT_0E (INIT_0E),
               .INIT_0F (INIT_0F),
               .INIT_10 (INIT_10),
               .INIT_11 (INIT_11),
               .INIT_12 (INIT_12),
               .INIT_13 (INIT_13),
               .INIT_14 (INIT_14),
               .INIT_15 (INIT_15),
               .INIT_16 (INIT_16),
               .INIT_17 (INIT_17),
               .INIT_18 (INIT_18),
               .INIT_19 (INIT_19),
               .INIT_1A (INIT_1A),
               .INIT_1B (INIT_1B),
               .INIT_1C (INIT_1C),
               .INIT_1D (INIT_1D),
               .INIT_1E (INIT_1E),
               .INIT_1F (INIT_1F),
               .INIT_20 (INIT_20),
               .INIT_21 (INIT_21),
               .INIT_22 (INIT_22),
               .INIT_23 (INIT_23),
               .INIT_24 (INIT_24),
               .INIT_25 (INIT_25),
               .INIT_26 (INIT_26),
               .INIT_27 (INIT_27),
               .INIT_28 (INIT_28),
               .INIT_29 (INIT_29),
               .INIT_2A (INIT_2A),
               .INIT_2B (INIT_2B),
               .INIT_2C (INIT_2C),
               .INIT_2D (INIT_2D),
               .INIT_2E (INIT_2E),
               .INIT_2F (INIT_2F),
               .INIT_30 (INIT_30),
               .INIT_31 (INIT_31),
               .INIT_32 (INIT_32),
               .INIT_33 (INIT_33),
               .INIT_34 (INIT_34),
               .INIT_35 (INIT_35),
               .INIT_36 (INIT_36),
               .INIT_37 (INIT_37),
               .INIT_38 (INIT_38),
               .INIT_39 (INIT_39),
               .INIT_3A (INIT_3A),
               .INIT_3B (INIT_3B),
               .INIT_3C (INIT_3C),
               .INIT_3D (INIT_3D),
               .INIT_3E (INIT_3E),
               .INIT_3F (INIT_3F),
               .INIT_40 (INIT_40), 
               .INIT_41 (INIT_41),
               .INIT_42 (INIT_42),
               .INIT_43 (INIT_43),
               .INIT_44 (INIT_44),
               .INIT_45 (INIT_45),
               .INIT_46 (INIT_46),
               .INIT_47 (INIT_47),
               .INIT_48 (INIT_48),
               .INIT_49 (INIT_49),
               .INIT_4A (INIT_4A),
               .INIT_4B (INIT_4B),
               .INIT_4C (INIT_4C),
               .INIT_4D (INIT_4D),
               .INIT_4E (INIT_4E),
               .INIT_4F (INIT_4F),
               .INIT_50 (INIT_50),
               .INIT_51 (INIT_51),
               .INIT_52 (INIT_52),
               .INIT_53 (INIT_53),
               .INIT_54 (INIT_54),
               .INIT_55 (INIT_55),
               .INIT_56 (INIT_56),
               .INIT_57 (INIT_57),
               .INIT_58 (INIT_58),
               .INIT_59 (INIT_59),
               .INIT_5A (INIT_5A),
               .INIT_5B (INIT_5B),
               .INIT_5C (INIT_5C),
               .INIT_5D (INIT_5D),
               .INIT_5E (INIT_5E),
               .INIT_5F (INIT_5F),
               .INIT_60 (INIT_60),
               .INIT_61 (INIT_61),
               .INIT_62 (INIT_62),
               .INIT_63 (INIT_63),
               .INIT_64 (INIT_64),
               .INIT_65 (INIT_65),
               .INIT_66 (INIT_66),
               .INIT_67 (INIT_67),
               .INIT_68 (INIT_68),
               .INIT_69 (INIT_69),
               .INIT_6A (INIT_6A),
               .INIT_6B (INIT_6B),
               .INIT_6C (INIT_6C),
               .INIT_6D (INIT_6D),
               .INIT_6E (INIT_6E),
               .INIT_6F (INIT_6F),
               .INIT_70 (INIT_70),
               .INIT_71 (INIT_71),
               .INIT_72 (INIT_72),
               .INIT_73 (INIT_73),
               .INIT_74 (INIT_74),
               .INIT_75 (INIT_75),
               .INIT_76 (INIT_76),
               .INIT_77 (INIT_77),
               .INIT_78 (INIT_78),
               .INIT_79 (INIT_79),
               .INIT_7A (INIT_7A),
               .INIT_7B (INIT_7B),
               .INIT_7C (INIT_7C),
               .INIT_7D (INIT_7D),
               .INIT_7E (INIT_7E),
               .INIT_7F (INIT_7F),
               .INIT_FILE (INIT_FILE),
               .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
               .SIM_MODE (SIM_MODE),
               .SRVAL(srval_tmp) 
               ) bram36_sdp (
               .DBITERR (),
               .DO (DO_PATTERN), 
               .DOP (DOP_PATTERN), 
               .ECCPARITY(), 
               .SBITERR (),
               .DI (DI_PATTERN), 
               .DIP (DIP_PATTERN), 
               .RDADDR (RDADDR), 
               .RDCLK (RDCLK), 
               .RDEN (RDEN), 
               .REGCE (REGCE), 
               .SSR (RST),  
               .WE (WE_PATTERN), 
               .WRADDR (WRADDR), 
               .WRCLK (WRCLK), 
               .WREN (WREN)
               );
             end 
           end // end generate virtex5
          // begin generate virtex6
         "VIRTEX6", "7SERIES" : 
           begin
             if (BRAM_SIZE == "18Kb" && READ_WIDTH <= 18 && WRITE_WIDTH <= 18) begin : bram18_dp_bl
              RAMB18E1 # ( 
                .DOA_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A (init_tmp),
                .INIT_B (init_tmp),
                .INIT_FILE(INIT_FILE),
                .RAM_MODE("TDP"),
                .READ_WIDTH_A (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_DEVICE ("7SERIES"),
                .SRVAL_A (srval_tmp),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE),
                .WRITE_WIDTH_B (wr_width)
                )  bram18_tdp_bl (
                .DOADO (DO_PATTERN[15:0]), 
                .DOBDO (), 
                .DOPADOP (DOP_PATTERN[1:0]), 
                .DOPBDOP (),
                .ADDRARDADDR (RDADDR_PATTERN), 
                .ADDRBWRADDR (WRADDR_PATTERN), 
                .CLKARDCLK (RDCLK), 
                .CLKBWRCLK (WRCLK), 
                .DIADI (16'b0), 
                .DIBDI (DI_PATTERN[15:0]), 
                .DIPADIP (2'b0), 
                .DIPBDIP (DIP_PATTERN[1:0]), 
                .ENARDEN (RDEN), 
                .ENBWREN (WREN), 
                .REGCEAREGCE (REGCE), 
                .REGCEB (1'b0), 
                .RSTRAMARSTRAM (RSTRAM_PATTERN), 
                .RSTRAMB (RSTRAM_PATTERN), 
                .RSTREGARSTREG (RSTREG_PATTERN), 
                .RSTREGB (RSTREG_PATTERN), 
                .WEA (2'b0), 
                .WEBWE (WE_PATTERN)
                );
              end
             else if (BRAM_SIZE == "18Kb" && ( (READ_WIDTH > 18 && READ_WIDTH <= 36) && (WRITE_WIDTH <= 18)) ) begin : bram18_sdp_bl_1
               RAMB18E1 # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A ({init_tmp[33:32],init_tmp[15:0]}),
                .INIT_B ({init_tmp[35:34],init_tmp[31:16]}),
                .INIT_FILE(INIT_FILE),
                .RAM_MODE("SDP"),
                .READ_WIDTH_A (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_DEVICE ("7SERIES"),
                .SRVAL_A ({srval_tmp[33:32],srval_tmp[15:0]}),
                .SRVAL_B ({srval_tmp[35:34],srval_tmp[31:16]}),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE),
                .WRITE_WIDTH_B (wr_width)
                )  bram18_sdp_bl_1 (
                .DOADO (DO_PATTERN[15:0]), 
                .DOBDO (DO_PATTERN[31:16]), 
                .DOPADOP (DOP_PATTERN[1:0]),
                .DOPBDOP (DOP_PATTERN[3:2]), 
                .ADDRARDADDR (RDADDR_PATTERN), 
                .ADDRBWRADDR (WRADDR_PATTERN), 
                .CLKARDCLK (RDCLK), 
                .CLKBWRCLK (WRCLK), 
                .DIADI (16'b0), 
                .DIBDI (DI_PATTERN[15:0]), 
                .DIPADIP (2'b0), 
                .DIPBDIP (DIP_PATTERN[1:0]), 
                .ENARDEN (RDEN), 
                .ENBWREN (WREN), 
                .REGCEAREGCE (REGCE), 
                .REGCEB (1'b0), 
                .RSTRAMARSTRAM (RSTRAM_PATTERN), 
                .RSTRAMB (RSTRAM_PATTERN), 
                .RSTREGARSTREG (RSTREG_PATTERN), 
                .RSTREGB (RSTREG_PATTERN), 
                .WEA (2'b0), 
                .WEBWE (WE_PATTERN)
                );
              end 
          else if (BRAM_SIZE == "18Kb" && ( (READ_WIDTH <= 18) && (WRITE_WIDTH > 18  && WRITE_WIDTH <= 36)) ) begin : bram18_sdp_bl_2
               RAMB18E1 # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A ({init_tmp[33:32],init_tmp[15:0]}),
                .INIT_B ({init_tmp[35:34],init_tmp[31:16]}),
                .INIT_FILE(INIT_FILE),
                .RAM_MODE("SDP"),
                .READ_WIDTH_A (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_DEVICE ("7SERIES"),
                .SRVAL_A ({srval_tmp[33:32],srval_tmp[15:0]}),
                .SRVAL_B ({srval_tmp[35:34],srval_tmp[31:16]}),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE),
                .WRITE_WIDTH_B (wr_width)
                )  bram18_sdp_bl_1 (
                .DOADO (DO_PATTERN[15:0]), 
                .DOBDO (), 
                .DOPADOP (DOP_PATTERN[1:0]),
                .DOPBDOP (), 
                .ADDRARDADDR (RDADDR_PATTERN), 
                .ADDRBWRADDR (WRADDR_PATTERN), 
                .CLKARDCLK (RDCLK), 
                .CLKBWRCLK (WRCLK), 
                .DIADI (DI_PATTERN[15:0]), 
                .DIBDI (DI_PATTERN[31:16]), 
                .DIPADIP (DIP_PATTERN[1:0]), 
                .DIPBDIP (DIP_PATTERN[3:2]), 
                .ENARDEN (RDEN), 
                .ENBWREN (WREN), 
                .REGCEAREGCE (REGCE), 
                .REGCEB (1'b0), 
                .RSTRAMARSTRAM (RSTRAM_PATTERN), 
                .RSTRAMB (RSTRAM_PATTERN), 
                .RSTREGARSTREG (RSTREG_PATTERN), 
                .RSTREGB (RSTREG_PATTERN), 
                .WEA (2'b0), 
                .WEBWE (WE_PATTERN)
                );
              end 
           else if (BRAM_SIZE == "18Kb" && ( (READ_WIDTH > 18 && READ_WIDTH <= 36) && (WRITE_WIDTH > 18  && WRITE_WIDTH <= 36)) ) begin : bram18_sdp_bl_3
               RAMB18E1 # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A ({init_tmp[33:32],init_tmp[15:0]}),
                .INIT_B ({init_tmp[35:34],init_tmp[31:16]}),
                .INIT_FILE(INIT_FILE),
                .RAM_MODE("SDP"),
                .READ_WIDTH_A (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_DEVICE ("7SERIES"),
                .SRVAL_A ({srval_tmp[33:32],srval_tmp[15:0]}),
                .SRVAL_B ({srval_tmp[35:34],srval_tmp[31:16]}),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE),
                .WRITE_WIDTH_B (wr_width)
                )  bram18_sdp_bl_3 (
                .DOADO (DO_PATTERN[15:0]), 
                .DOBDO (DO_PATTERN[31:16]), 
                .DOPADOP (DOP_PATTERN[1:0]),
                .DOPBDOP (DOP_PATTERN[3:2]), 
                .ADDRARDADDR (RDADDR_PATTERN), 
                .ADDRBWRADDR (WRADDR_PATTERN), 
                .CLKARDCLK (RDCLK), 
                .CLKBWRCLK (WRCLK), 
                .DIADI (DI_PATTERN[15:0]), 
                .DIBDI (DI_PATTERN[31:16]), 
                .DIPADIP (DIP_PATTERN[1:0]), 
                .DIPBDIP (DIP_PATTERN[3:2]), 
                .ENARDEN (RDEN), 
                .ENBWREN (WREN), 
                .REGCEAREGCE (REGCE), 
                .REGCEB (1'b0), 
                .RSTRAMARSTRAM (RSTRAM_PATTERN), 
                .RSTRAMB (RSTRAM_PATTERN), 
                .RSTREGARSTREG (RSTREG_PATTERN), 
                .RSTREGB (RSTREG_PATTERN), 
                .WEA (2'b0), 
                .WEBWE (WE_PATTERN)
                );
              end 
          else if (BRAM_SIZE == "36Kb" && (READ_WIDTH <= 36 && WRITE_WIDTH <= 36) ) begin : bram36_dp_bl
   
          RAMB36E1 # ( 
              .DOA_REG (DO_REG),
              .INITP_00 (INITP_00),
              .INITP_01 (INITP_01),
              .INITP_02 (INITP_02), 
              .INITP_03 (INITP_03),
              .INITP_04 (INITP_04),
              .INITP_05 (INITP_05),
              .INITP_06 (INITP_06),
              .INITP_07 (INITP_07),
	      .INITP_08 (INITP_08),
              .INITP_09 (INITP_09),
              .INITP_0A (INITP_0A),
              .INITP_0B (INITP_0B),
              .INITP_0C (INITP_0C),
              .INITP_0D (INITP_0D),
              .INITP_0E (INITP_0E),
              .INITP_0F (INITP_0F),
              .INIT_00 (INIT_00), 
              .INIT_01 (INIT_01),
              .INIT_02 (INIT_02),
              .INIT_03 (INIT_03),
              .INIT_04 (INIT_04),
              .INIT_05 (INIT_05),
              .INIT_06 (INIT_06),
              .INIT_07 (INIT_07),
              .INIT_08 (INIT_08),
              .INIT_09 (INIT_09),
              .INIT_0A (INIT_0A),
              .INIT_0B (INIT_0B),
              .INIT_0C (INIT_0C),
              .INIT_0D (INIT_0D),
              .INIT_0E (INIT_0E),
              .INIT_0F (INIT_0F),
              .INIT_10 (INIT_10),
              .INIT_11 (INIT_11),
              .INIT_12 (INIT_12),
              .INIT_13 (INIT_13),
              .INIT_14 (INIT_14),
              .INIT_15 (INIT_15),
              .INIT_16 (INIT_16),
              .INIT_17 (INIT_17),
              .INIT_18 (INIT_18),
              .INIT_19 (INIT_19),
              .INIT_1A (INIT_1A),
              .INIT_1B (INIT_1B),
              .INIT_1C (INIT_1C),
              .INIT_1D (INIT_1D),
              .INIT_1E (INIT_1E),
              .INIT_1F (INIT_1F),
              .INIT_20 (INIT_20),
              .INIT_21 (INIT_21),
              .INIT_22 (INIT_22),
              .INIT_23 (INIT_23),
              .INIT_24 (INIT_24),
              .INIT_25 (INIT_25),
              .INIT_26 (INIT_26),
              .INIT_27 (INIT_27),
              .INIT_28 (INIT_28),
              .INIT_29 (INIT_29),
              .INIT_2A (INIT_2A),
              .INIT_2B (INIT_2B),
              .INIT_2C (INIT_2C),
              .INIT_2D (INIT_2D),
              .INIT_2E (INIT_2E),
              .INIT_2F (INIT_2F),
              .INIT_30 (INIT_30),
              .INIT_31 (INIT_31),
              .INIT_32 (INIT_32),
              .INIT_33 (INIT_33),
              .INIT_34 (INIT_34),
              .INIT_35 (INIT_35),
              .INIT_36 (INIT_36),
              .INIT_37 (INIT_37),
              .INIT_38 (INIT_38),
              .INIT_39 (INIT_39),
              .INIT_3A (INIT_3A),
              .INIT_3B (INIT_3B),
              .INIT_3C (INIT_3C),
              .INIT_3D (INIT_3D),
              .INIT_3E (INIT_3E),
              .INIT_3F (INIT_3F),
              .INIT_40 (INIT_40), 
              .INIT_41 (INIT_41),
              .INIT_42 (INIT_42),
              .INIT_43 (INIT_43),
              .INIT_44 (INIT_44),
              .INIT_45 (INIT_45),
              .INIT_46 (INIT_46),
              .INIT_47 (INIT_47),
              .INIT_48 (INIT_48),
              .INIT_49 (INIT_49),
              .INIT_4A (INIT_4A),
              .INIT_4B (INIT_4B),
              .INIT_4C (INIT_4C),
              .INIT_4D (INIT_4D),
              .INIT_4E (INIT_4E),
              .INIT_4F (INIT_4F),
              .INIT_50 (INIT_50),
              .INIT_51 (INIT_51),
              .INIT_52 (INIT_52),
              .INIT_53 (INIT_53),
              .INIT_54 (INIT_54),
              .INIT_55 (INIT_55),
              .INIT_56 (INIT_56),
              .INIT_57 (INIT_57),
              .INIT_58 (INIT_58),
              .INIT_59 (INIT_59),
              .INIT_5A (INIT_5A),
              .INIT_5B (INIT_5B),
              .INIT_5C (INIT_5C),
              .INIT_5D (INIT_5D),
              .INIT_5E (INIT_5E),
              .INIT_5F (INIT_5F),
              .INIT_60 (INIT_60),
              .INIT_61 (INIT_61),
              .INIT_62 (INIT_62),
              .INIT_63 (INIT_63),
              .INIT_64 (INIT_64),
              .INIT_65 (INIT_65),
              .INIT_66 (INIT_66),
              .INIT_67 (INIT_67),
              .INIT_68 (INIT_68),
              .INIT_69 (INIT_69),
              .INIT_6A (INIT_6A),
              .INIT_6B (INIT_6B),
              .INIT_6C (INIT_6C),
              .INIT_6D (INIT_6D),
              .INIT_6E (INIT_6E),
              .INIT_6F (INIT_6F),
              .INIT_70 (INIT_70),
              .INIT_71 (INIT_71),
              .INIT_72 (INIT_72),
              .INIT_73 (INIT_73),
              .INIT_74 (INIT_74),
              .INIT_75 (INIT_75),
              .INIT_76 (INIT_76),
              .INIT_77 (INIT_77),
              .INIT_78 (INIT_78),
              .INIT_79 (INIT_79),
              .INIT_7A (INIT_7A),
              .INIT_7B (INIT_7B),
              .INIT_7C (INIT_7C),
              .INIT_7D (INIT_7D),
              .INIT_7E (INIT_7E),
              .INIT_7F (INIT_7F),
              .INIT_A (init_tmp),
              .INIT_FILE (INIT_FILE),
              .RAM_MODE ("TDP"),
              .READ_WIDTH_A (rd_width),
              .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
              .SIM_DEVICE ("7SERIES"),
              .SRVAL_A (srval_tmp),
              .WRITE_MODE_A (WRITE_MODE),
              .WRITE_MODE_B (WRITE_MODE),
              .WRITE_WIDTH_B (wr_width)
              )  bram36_tdp_bl (
              .CASCADEOUTA (),
              .CASCADEOUTB (),
              .DBITERR (),
              .DOADO (DO_PATTERN), 
              .DOBDO (), 
              .DOPADOP (DOP_PATTERN), 
              .DOPBDOP (),
              .ECCPARITY (),
              .RDADDRECC (),
              .SBITERR (),
              .ADDRARDADDR (RDADDR_PATTERN), 
              .ADDRBWRADDR (WRADDR_PATTERN),
              .CASCADEINA (1'b0),
              .CASCADEINB (1'b0), 
              .CLKARDCLK (RDCLK), 
              .CLKBWRCLK (WRCLK), 
              .DIADI (32'b0), 
              .DIBDI (DI_PATTERN), 
              .DIPADIP (4'b0), 
              .DIPBDIP (DIP_PATTERN), 
              .ENARDEN (RDEN), 
              .ENBWREN (WREN), 
              .INJECTDBITERR(1'b0),
              .INJECTSBITERR(1'b0),
              .REGCEAREGCE (REGCE), 
              .REGCEB (1'b0), 
              .RSTRAMARSTRAM (RSTRAM_PATTERN), 
              .RSTRAMB (RSTRAM_PATTERN), 
              .RSTREGARSTREG (RSTREG_PATTERN), 
              .RSTREGB (RSTREG_PATTERN), 
              .WEA (4'b0), 
              .WEBWE (WE_PATTERN)
              );
            end

            else if (BRAM_SIZE == "36Kb" && ( (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) && (READ_WIDTH <= 36) ) ) begin : bram36_sdp_bl
   
            RAMB36E1 # ( 
              .DOA_REG (DO_REG),
              .DOB_REG (DO_REG),
              .INITP_00 (INITP_00),
              .INITP_01 (INITP_01),
              .INITP_02 (INITP_02), 
              .INITP_03 (INITP_03),
              .INITP_04 (INITP_04),
              .INITP_05 (INITP_05),
              .INITP_06 (INITP_06),
              .INITP_07 (INITP_07),
	      .INITP_08 (INITP_08),
              .INITP_09 (INITP_09),
              .INITP_0A (INITP_0A),
              .INITP_0B (INITP_0B),
              .INITP_0C (INITP_0C),
              .INITP_0D (INITP_0D),
              .INITP_0E (INITP_0E),
              .INITP_0F (INITP_0F),
              .INIT_00 (INIT_00), 
              .INIT_01 (INIT_01),
              .INIT_02 (INIT_02),
              .INIT_03 (INIT_03),
              .INIT_04 (INIT_04),
              .INIT_05 (INIT_05),
              .INIT_06 (INIT_06),
              .INIT_07 (INIT_07),
              .INIT_08 (INIT_08),
              .INIT_09 (INIT_09),
              .INIT_0A (INIT_0A),
              .INIT_0B (INIT_0B),
              .INIT_0C (INIT_0C),
              .INIT_0D (INIT_0D),
              .INIT_0E (INIT_0E),
              .INIT_0F (INIT_0F),
              .INIT_10 (INIT_10),
              .INIT_11 (INIT_11),
              .INIT_12 (INIT_12),
              .INIT_13 (INIT_13),
              .INIT_14 (INIT_14),
              .INIT_15 (INIT_15),
              .INIT_16 (INIT_16),
              .INIT_17 (INIT_17),
              .INIT_18 (INIT_18),
              .INIT_19 (INIT_19),
              .INIT_1A (INIT_1A),
              .INIT_1B (INIT_1B),
              .INIT_1C (INIT_1C),
              .INIT_1D (INIT_1D),
              .INIT_1E (INIT_1E),
              .INIT_1F (INIT_1F),
              .INIT_20 (INIT_20),
              .INIT_21 (INIT_21),
              .INIT_22 (INIT_22),
              .INIT_23 (INIT_23),
              .INIT_24 (INIT_24),
              .INIT_25 (INIT_25),
              .INIT_26 (INIT_26),
              .INIT_27 (INIT_27),
              .INIT_28 (INIT_28),
              .INIT_29 (INIT_29),
              .INIT_2A (INIT_2A),
              .INIT_2B (INIT_2B),
              .INIT_2C (INIT_2C),
              .INIT_2D (INIT_2D),
              .INIT_2E (INIT_2E),
              .INIT_2F (INIT_2F),
              .INIT_30 (INIT_30),
              .INIT_31 (INIT_31),
              .INIT_32 (INIT_32),
              .INIT_33 (INIT_33),
              .INIT_34 (INIT_34),
              .INIT_35 (INIT_35),
              .INIT_36 (INIT_36),
              .INIT_37 (INIT_37),
              .INIT_38 (INIT_38),
              .INIT_39 (INIT_39),
              .INIT_3A (INIT_3A),
              .INIT_3B (INIT_3B),
              .INIT_3C (INIT_3C),
              .INIT_3D (INIT_3D),
              .INIT_3E (INIT_3E),
              .INIT_3F (INIT_3F),
              .INIT_40 (INIT_40), 
              .INIT_41 (INIT_41),
              .INIT_42 (INIT_42),
              .INIT_43 (INIT_43),
              .INIT_44 (INIT_44),
              .INIT_45 (INIT_45),
              .INIT_46 (INIT_46),
              .INIT_47 (INIT_47),
              .INIT_48 (INIT_48),
              .INIT_49 (INIT_49),
              .INIT_4A (INIT_4A),
              .INIT_4B (INIT_4B),
              .INIT_4C (INIT_4C),
              .INIT_4D (INIT_4D),
              .INIT_4E (INIT_4E),
              .INIT_4F (INIT_4F),
              .INIT_50 (INIT_50),
              .INIT_51 (INIT_51),
              .INIT_52 (INIT_52),
              .INIT_53 (INIT_53),
              .INIT_54 (INIT_54),
              .INIT_55 (INIT_55),
              .INIT_56 (INIT_56),
              .INIT_57 (INIT_57),
              .INIT_58 (INIT_58),
              .INIT_59 (INIT_59),
              .INIT_5A (INIT_5A),
              .INIT_5B (INIT_5B),
              .INIT_5C (INIT_5C),
              .INIT_5D (INIT_5D),
              .INIT_5E (INIT_5E),
              .INIT_5F (INIT_5F),
              .INIT_60 (INIT_60),
              .INIT_61 (INIT_61),
              .INIT_62 (INIT_62),
              .INIT_63 (INIT_63),
              .INIT_64 (INIT_64),
              .INIT_65 (INIT_65),
              .INIT_66 (INIT_66),
              .INIT_67 (INIT_67),
              .INIT_68 (INIT_68),
              .INIT_69 (INIT_69),
              .INIT_6A (INIT_6A),
              .INIT_6B (INIT_6B),
              .INIT_6C (INIT_6C),
              .INIT_6D (INIT_6D),
              .INIT_6E (INIT_6E),
              .INIT_6F (INIT_6F),
              .INIT_70 (INIT_70),
              .INIT_71 (INIT_71),
              .INIT_72 (INIT_72),
              .INIT_73 (INIT_73),
              .INIT_74 (INIT_74),
              .INIT_75 (INIT_75),
              .INIT_76 (INIT_76),
              .INIT_77 (INIT_77),
              .INIT_78 (INIT_78),
              .INIT_79 (INIT_79),
              .INIT_7A (INIT_7A),
              .INIT_7B (INIT_7B),
              .INIT_7C (INIT_7C),
              .INIT_7D (INIT_7D),
              .INIT_7E (INIT_7E),
              .INIT_7F (INIT_7F),
              .INIT_A ({init_tmp[67:64],init_tmp[31:0]}),
              .INIT_B ({init_tmp[71:68],init_tmp[63:32]}),
              .INIT_FILE (INIT_FILE),
              .RAM_MODE ("SDP"),
              .READ_WIDTH_A (rd_width),
              .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
              .SIM_DEVICE ("7SERIES"),
              .SRVAL_A ({srval_tmp[67:64],srval_tmp[31:0]}),
              .SRVAL_B ({srval_tmp[71:68],srval_tmp[63:32]}),
              .WRITE_MODE_A (WRITE_MODE),
              .WRITE_MODE_B (WRITE_MODE),
              .WRITE_WIDTH_B (wr_width)
              )  bram36_sdp_bl (
              .CASCADEOUTA (),
              .CASCADEOUTB (),
              .DBITERR (),
              .DOADO (DO_PATTERN[31:0]), 
              .DOBDO (), 
              .DOPADOP (DOP_PATTERN[3:0]), 
              .DOPBDOP (),
              .ECCPARITY (),
              .RDADDRECC (),
              .SBITERR (),
              .ADDRARDADDR (RDADDR_PATTERN), 
              .ADDRBWRADDR (WRADDR_PATTERN),
              .CASCADEINA (1'b0),
              .CASCADEINB (1'b0), 
              .CLKARDCLK (RDCLK), 
              .CLKBWRCLK (WRCLK), 
              .DIADI (DI_PATTERN[31:0]), 
              .DIBDI (DI_PATTERN[63:32]), 
              .DIPADIP (DIP_PATTERN[3:0]), 
              .DIPBDIP (DIP_PATTERN[7:4]), 
              .ENARDEN (RDEN), 
              .ENBWREN (WREN), 
              .INJECTDBITERR(1'b0),
              .INJECTSBITERR(1'b0),
              .REGCEAREGCE (REGCE), 
              .REGCEB (1'b0), 
              .RSTRAMARSTRAM (RSTRAM_PATTERN), 
              .RSTRAMB (RSTRAM_PATTERN), 
              .RSTREGARSTREG (RSTREG_PATTERN), 
              .RSTREGB (RSTREG_PATTERN), 
              .WEA (4'b0), 
              .WEBWE (WE_PATTERN)
              );
            
             end 
             else if (BRAM_SIZE == "36Kb" && ( (READ_WIDTH > 36 && READ_WIDTH <= 72) && (WRITE_WIDTH <= 36) ) ) begin : bram36_sdp_bl_1
   
            RAMB36E1 # ( 
              .DOA_REG (DO_REG),
              .DOB_REG (DO_REG),
              .INITP_00 (INITP_00),
              .INITP_01 (INITP_01),
              .INITP_02 (INITP_02), 
              .INITP_03 (INITP_03),
              .INITP_04 (INITP_04),
              .INITP_05 (INITP_05),
              .INITP_06 (INITP_06),
              .INITP_07 (INITP_07),
	      .INITP_08 (INITP_08),
              .INITP_09 (INITP_09),
              .INITP_0A (INITP_0A),
              .INITP_0B (INITP_0B),
              .INITP_0C (INITP_0C),
              .INITP_0D (INITP_0D),
              .INITP_0E (INITP_0E),
              .INITP_0F (INITP_0F),			 
              .INIT_00 (INIT_00), 
              .INIT_01 (INIT_01),
              .INIT_02 (INIT_02),
              .INIT_03 (INIT_03),
              .INIT_04 (INIT_04),
              .INIT_05 (INIT_05),
              .INIT_06 (INIT_06),
              .INIT_07 (INIT_07),
              .INIT_08 (INIT_08),
              .INIT_09 (INIT_09),
              .INIT_0A (INIT_0A),
              .INIT_0B (INIT_0B),
              .INIT_0C (INIT_0C),
              .INIT_0D (INIT_0D),
              .INIT_0E (INIT_0E),
              .INIT_0F (INIT_0F),
              .INIT_10 (INIT_10),
              .INIT_11 (INIT_11),
              .INIT_12 (INIT_12),
              .INIT_13 (INIT_13),
              .INIT_14 (INIT_14),
              .INIT_15 (INIT_15),
              .INIT_16 (INIT_16),
              .INIT_17 (INIT_17),
              .INIT_18 (INIT_18),
              .INIT_19 (INIT_19),
              .INIT_1A (INIT_1A),
              .INIT_1B (INIT_1B),
              .INIT_1C (INIT_1C),
              .INIT_1D (INIT_1D),
              .INIT_1E (INIT_1E),
              .INIT_1F (INIT_1F),
              .INIT_20 (INIT_20),
              .INIT_21 (INIT_21),
              .INIT_22 (INIT_22),
              .INIT_23 (INIT_23),
              .INIT_24 (INIT_24),
              .INIT_25 (INIT_25),
              .INIT_26 (INIT_26),
              .INIT_27 (INIT_27),
              .INIT_28 (INIT_28),
              .INIT_29 (INIT_29),
              .INIT_2A (INIT_2A),
              .INIT_2B (INIT_2B),
              .INIT_2C (INIT_2C),
              .INIT_2D (INIT_2D),
              .INIT_2E (INIT_2E),
              .INIT_2F (INIT_2F),
              .INIT_30 (INIT_30),
              .INIT_31 (INIT_31),
              .INIT_32 (INIT_32),
              .INIT_33 (INIT_33),
              .INIT_34 (INIT_34),
              .INIT_35 (INIT_35),
              .INIT_36 (INIT_36),
              .INIT_37 (INIT_37),
              .INIT_38 (INIT_38),
              .INIT_39 (INIT_39),
              .INIT_3A (INIT_3A),
              .INIT_3B (INIT_3B),
              .INIT_3C (INIT_3C),
              .INIT_3D (INIT_3D),
              .INIT_3E (INIT_3E),
              .INIT_3F (INIT_3F),
              .INIT_40 (INIT_40), 
              .INIT_41 (INIT_41),
              .INIT_42 (INIT_42),
              .INIT_43 (INIT_43),
              .INIT_44 (INIT_44),
              .INIT_45 (INIT_45),
              .INIT_46 (INIT_46),
              .INIT_47 (INIT_47),
              .INIT_48 (INIT_48),
              .INIT_49 (INIT_49),
              .INIT_4A (INIT_4A),
              .INIT_4B (INIT_4B),
              .INIT_4C (INIT_4C),
              .INIT_4D (INIT_4D),
              .INIT_4E (INIT_4E),
              .INIT_4F (INIT_4F),
              .INIT_50 (INIT_50),
              .INIT_51 (INIT_51),
              .INIT_52 (INIT_52),
              .INIT_53 (INIT_53),
              .INIT_54 (INIT_54),
              .INIT_55 (INIT_55),
              .INIT_56 (INIT_56),
              .INIT_57 (INIT_57),
              .INIT_58 (INIT_58),
              .INIT_59 (INIT_59),
              .INIT_5A (INIT_5A),
              .INIT_5B (INIT_5B),
              .INIT_5C (INIT_5C),
              .INIT_5D (INIT_5D),
              .INIT_5E (INIT_5E),
              .INIT_5F (INIT_5F),
              .INIT_60 (INIT_60),
              .INIT_61 (INIT_61),
              .INIT_62 (INIT_62),
              .INIT_63 (INIT_63),
              .INIT_64 (INIT_64),
              .INIT_65 (INIT_65),
              .INIT_66 (INIT_66),
              .INIT_67 (INIT_67),
              .INIT_68 (INIT_68),
              .INIT_69 (INIT_69),
              .INIT_6A (INIT_6A),
              .INIT_6B (INIT_6B),
              .INIT_6C (INIT_6C),
              .INIT_6D (INIT_6D),
              .INIT_6E (INIT_6E),
              .INIT_6F (INIT_6F),
              .INIT_70 (INIT_70),
              .INIT_71 (INIT_71),
              .INIT_72 (INIT_72),
              .INIT_73 (INIT_73),
              .INIT_74 (INIT_74),
              .INIT_75 (INIT_75),
              .INIT_76 (INIT_76),
              .INIT_77 (INIT_77),
              .INIT_78 (INIT_78),
              .INIT_79 (INIT_79),
              .INIT_7A (INIT_7A),
              .INIT_7B (INIT_7B),
              .INIT_7C (INIT_7C),
              .INIT_7D (INIT_7D),
              .INIT_7E (INIT_7E),
              .INIT_7F (INIT_7F),
              .INIT_A ({init_tmp[67:64],init_tmp[31:0]}),
              .INIT_B ({init_tmp[71:68],init_tmp[63:32]}),
              .INIT_FILE (INIT_FILE),
              .RAM_MODE ("SDP"),
              .READ_WIDTH_A (rd_width),
              .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
              .SIM_DEVICE ("7SERIES"),
              .SRVAL_A ({srval_tmp[67:64],srval_tmp[31:0]}),
              .SRVAL_B ({srval_tmp[71:68],srval_tmp[63:32]}),
              .WRITE_MODE_A (WRITE_MODE),
              .WRITE_MODE_B (WRITE_MODE),
              .WRITE_WIDTH_B (wr_width)
              )  bram36_sdp_bl_1 (
              .CASCADEOUTA (),
              .CASCADEOUTB (),
              .DBITERR (),
              .DOADO (DO_PATTERN[31:0]), 
              .DOBDO (DO_PATTERN[63:32]), 
              .DOPADOP (DOP_PATTERN[3:0]), 
              .DOPBDOP (DOP_PATTERN[7:4]),
              .ECCPARITY (),
              .RDADDRECC (),
              .SBITERR (),
              .ADDRARDADDR (RDADDR_PATTERN), 
              .ADDRBWRADDR (WRADDR_PATTERN),
              .CASCADEINA (1'b0),
              .CASCADEINB (1'b0), 
              .CLKARDCLK (RDCLK), 
              .CLKBWRCLK (WRCLK), 
              .DIADI (32'b0), 
              .DIBDI (DI_PATTERN[31:0]), 
              .DIPADIP (4'b0), 
              .DIPBDIP (DIP_PATTERN[3:0]), 
              .ENARDEN (RDEN), 
              .ENBWREN (WREN), 
              .INJECTDBITERR(1'b0),
              .INJECTSBITERR(1'b0),
              .REGCEAREGCE (REGCE), 
              .REGCEB (1'b0), 
              .RSTRAMARSTRAM (RSTRAM_PATTERN), 
              .RSTRAMB (RSTRAM_PATTERN), 
              .RSTREGARSTREG (RSTREG_PATTERN), 
              .RSTREGB (RSTREG_PATTERN), 
              .WEA (4'b0), 
              .WEBWE (WE_PATTERN)
              );
            
             end 
            else if (BRAM_SIZE == "36Kb" && ( (READ_WIDTH > 36 && READ_WIDTH <= 72) && (WRITE_WIDTH > 36 && WRITE_WIDTH <= 72) ) ) begin : bram36_sdp_bl_2
   
            RAMB36E1 # ( 
              .DOA_REG (DO_REG),
              .DOB_REG (DO_REG),
              .INITP_00 (INITP_00),
              .INITP_01 (INITP_01),
              .INITP_02 (INITP_02), 
              .INITP_03 (INITP_03),
              .INITP_04 (INITP_04),
              .INITP_05 (INITP_05),
              .INITP_06 (INITP_06),
              .INITP_07 (INITP_07),
	      .INITP_08 (INITP_08),
              .INITP_09 (INITP_09),
              .INITP_0A (INITP_0A),
              .INITP_0B (INITP_0B),
              .INITP_0C (INITP_0C),
              .INITP_0D (INITP_0D),
              .INITP_0E (INITP_0E),
              .INITP_0F (INITP_0F),
              .INIT_00 (INIT_00), 
              .INIT_01 (INIT_01),
              .INIT_02 (INIT_02),
              .INIT_03 (INIT_03),
              .INIT_04 (INIT_04),
              .INIT_05 (INIT_05),
              .INIT_06 (INIT_06),
              .INIT_07 (INIT_07),
              .INIT_08 (INIT_08),
              .INIT_09 (INIT_09),
              .INIT_0A (INIT_0A),
              .INIT_0B (INIT_0B),
              .INIT_0C (INIT_0C),
              .INIT_0D (INIT_0D),
              .INIT_0E (INIT_0E),
              .INIT_0F (INIT_0F),
              .INIT_10 (INIT_10),
              .INIT_11 (INIT_11),
              .INIT_12 (INIT_12),
              .INIT_13 (INIT_13),
              .INIT_14 (INIT_14),
              .INIT_15 (INIT_15),
              .INIT_16 (INIT_16),
              .INIT_17 (INIT_17),
              .INIT_18 (INIT_18),
              .INIT_19 (INIT_19),
              .INIT_1A (INIT_1A),
              .INIT_1B (INIT_1B),
              .INIT_1C (INIT_1C),
              .INIT_1D (INIT_1D),
              .INIT_1E (INIT_1E),
              .INIT_1F (INIT_1F),
              .INIT_20 (INIT_20),
              .INIT_21 (INIT_21),
              .INIT_22 (INIT_22),
              .INIT_23 (INIT_23),
              .INIT_24 (INIT_24),
              .INIT_25 (INIT_25),
              .INIT_26 (INIT_26),
              .INIT_27 (INIT_27),
              .INIT_28 (INIT_28),
              .INIT_29 (INIT_29),
              .INIT_2A (INIT_2A),
              .INIT_2B (INIT_2B),
              .INIT_2C (INIT_2C),
              .INIT_2D (INIT_2D),
              .INIT_2E (INIT_2E),
              .INIT_2F (INIT_2F),
              .INIT_30 (INIT_30),
              .INIT_31 (INIT_31),
              .INIT_32 (INIT_32),
              .INIT_33 (INIT_33),
              .INIT_34 (INIT_34),
              .INIT_35 (INIT_35),
              .INIT_36 (INIT_36),
              .INIT_37 (INIT_37),
              .INIT_38 (INIT_38),
              .INIT_39 (INIT_39),
              .INIT_3A (INIT_3A),
              .INIT_3B (INIT_3B),
              .INIT_3C (INIT_3C),
              .INIT_3D (INIT_3D),
              .INIT_3E (INIT_3E),
              .INIT_3F (INIT_3F),
              .INIT_40 (INIT_40), 
              .INIT_41 (INIT_41),
              .INIT_42 (INIT_42),
              .INIT_43 (INIT_43),
              .INIT_44 (INIT_44),
              .INIT_45 (INIT_45),
              .INIT_46 (INIT_46),
              .INIT_47 (INIT_47),
              .INIT_48 (INIT_48),
              .INIT_49 (INIT_49),
              .INIT_4A (INIT_4A),
              .INIT_4B (INIT_4B),
              .INIT_4C (INIT_4C),
              .INIT_4D (INIT_4D),
              .INIT_4E (INIT_4E),
              .INIT_4F (INIT_4F),
              .INIT_50 (INIT_50),
              .INIT_51 (INIT_51),
              .INIT_52 (INIT_52),
              .INIT_53 (INIT_53),
              .INIT_54 (INIT_54),
              .INIT_55 (INIT_55),
              .INIT_56 (INIT_56),
              .INIT_57 (INIT_57),
              .INIT_58 (INIT_58),
              .INIT_59 (INIT_59),
              .INIT_5A (INIT_5A),
              .INIT_5B (INIT_5B),
              .INIT_5C (INIT_5C),
              .INIT_5D (INIT_5D),
              .INIT_5E (INIT_5E),
              .INIT_5F (INIT_5F),
              .INIT_60 (INIT_60),
              .INIT_61 (INIT_61),
              .INIT_62 (INIT_62),
              .INIT_63 (INIT_63),
              .INIT_64 (INIT_64),
              .INIT_65 (INIT_65),
              .INIT_66 (INIT_66),
              .INIT_67 (INIT_67),
              .INIT_68 (INIT_68),
              .INIT_69 (INIT_69),
              .INIT_6A (INIT_6A),
              .INIT_6B (INIT_6B),
              .INIT_6C (INIT_6C),
              .INIT_6D (INIT_6D),
              .INIT_6E (INIT_6E),
              .INIT_6F (INIT_6F),
              .INIT_70 (INIT_70),
              .INIT_71 (INIT_71),
              .INIT_72 (INIT_72),
              .INIT_73 (INIT_73),
              .INIT_74 (INIT_74),
              .INIT_75 (INIT_75),
              .INIT_76 (INIT_76),
              .INIT_77 (INIT_77),
              .INIT_78 (INIT_78),
              .INIT_79 (INIT_79),
              .INIT_7A (INIT_7A),
              .INIT_7B (INIT_7B),
              .INIT_7C (INIT_7C),
              .INIT_7D (INIT_7D),
              .INIT_7E (INIT_7E),
              .INIT_7F (INIT_7F),
              .INIT_A ({init_tmp[67:64],init_tmp[31:0]}),
              .INIT_B ({init_tmp[71:68],init_tmp[63:32]}),
              .INIT_FILE (INIT_FILE),
              .RAM_MODE ("SDP"),
              .READ_WIDTH_A (rd_width),
              .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
              .SIM_DEVICE ("7SERIES"),
              .SRVAL_A ({srval_tmp[67:64],srval_tmp[31:0]}),
              .SRVAL_B ({srval_tmp[71:68],srval_tmp[63:32]}),
              .WRITE_MODE_A (WRITE_MODE),
              .WRITE_MODE_B (WRITE_MODE),
              .WRITE_WIDTH_B (wr_width)
              )  bram36_sdp_bl_2 (
              .CASCADEOUTA (),
              .CASCADEOUTB (),
              .DBITERR (),
              .DOADO (DO_PATTERN[31:0]), 
              .DOBDO (DO_PATTERN[63:32]), 
              .DOPADOP (DOP_PATTERN[3:0]), 
              .DOPBDOP (DOP_PATTERN[7:4]),
              .ECCPARITY (),
              .RDADDRECC (),
              .SBITERR (),
              .ADDRARDADDR (RDADDR_PATTERN), 
              .ADDRBWRADDR (WRADDR_PATTERN),
              .CASCADEINA (1'b0),
              .CASCADEINB (1'b0), 
              .CLKARDCLK (RDCLK), 
              .CLKBWRCLK (WRCLK), 
              .DIADI (DI_PATTERN[31:0]), 
              .DIBDI (DI_PATTERN[63:32]), 
              .DIPADIP (DIP_PATTERN[3:0]), 
              .DIPBDIP (DIP_PATTERN[7:4]), 
              .ENARDEN (RDEN), 
              .ENBWREN (WREN), 
              .INJECTDBITERR(1'b0),
              .INJECTSBITERR(1'b0),
              .REGCEAREGCE (REGCE), 
              .REGCEB (1'b0), 
              .RSTRAMARSTRAM (RSTRAM_PATTERN), 
              .RSTRAMB (RSTRAM_PATTERN), 
              .RSTREGARSTREG (RSTREG_PATTERN), 
              .RSTREGB (RSTREG_PATTERN), 
              .WEA (4'b0), 
              .WEBWE (WE_PATTERN)
              );
            
             end 
           end  // end generate virtex6
       // begin generate spartan6
       "SPARTAN6" :  
          begin
            if (BRAM_SIZE == "9Kb" && WRITE_WIDTH <= 18) begin : bram9_tdp_stan
              RAMB8BWER # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_A (init_tmp),
                .INIT_B (init_tmp),
		.INIT_FILE (INIT_FILE),
                .DATA_WIDTH_A (wr_width),
                .DATA_WIDTH_B (rd_width),
                .RAM_MODE ("TDP"),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SRVAL_A (srval_tmp),
                .SRVAL_B (srval_tmp),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE)
                )  ram8bwe_tdp (
                .DOADO (), 
                .DOBDO (DO_PATTERN), 
                .DOPADOP (), 
                .DOPBDOP (DOP_PATTERN),
                .ADDRAWRADDR (WRADDR_PATTERN), 
                .ADDRBRDADDR (RDADDR_PATTERN), 
                .CLKAWRCLK (WRCLK), 
                .CLKBRDCLK (RDCLK), 
                .DIADI (DI_PATTERN), 
                .DIBDI (16'b0), 
                .DIPADIP (DIP_PATTERN), 
                .DIPBDIP (2'b0), 
                .ENAWREN (WREN), 
                .ENBRDEN (RDEN), 
                .REGCEA (1'b0), 
                .REGCEBREGCE (REGCE), 
                .RSTA (1'b0), 
                .RSTBRST (RST), 
                .WEAWEL (WE_PATTERN), 
                .WEBWEU (2'b0)
                );
            end
            else if (BRAM_SIZE == "9Kb" && WRITE_WIDTH > 18 && WRITE_WIDTH <= 36) begin : bram9_sdp_stan
              RAMB8BWER # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_A ({init_tmp[33:32],init_tmp[15:0]}),
                .INIT_B ({init_tmp[35:34],init_tmp[31:16]}),
		.INIT_FILE (INIT_FILE),
                .DATA_WIDTH_A (wr_width),
                .DATA_WIDTH_B (rd_width),
                .RAM_MODE ("SDP"),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SRVAL_A ({srval_tmp[33:32],srval_tmp[15:0]}),
                .SRVAL_B ({srval_tmp[35:34],srval_tmp[31:16]}),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE)
                )  ram8bwe_sdp (
                .DOADO (DO_PATTERN[15:0]), 
                .DOBDO (DO_PATTERN[31:16]), 
                .DOPADOP (DOP_PATTERN[1:0]), 
                .DOPBDOP (DOP_PATTERN[3:2]),
                .ADDRAWRADDR (WRADDR_PATTERN), 
                .ADDRBRDADDR (RDADDR_PATTERN), 
                .CLKAWRCLK (WRCLK), 
                .CLKBRDCLK (RDCLK), 
                .DIADI (DI_PATTERN[15:0]), 
                .DIBDI (DI_PATTERN[31:16]), 
                .DIPADIP (DIP_PATTERN[1:0]), 
                .DIPBDIP (DIP_PATTERN[3:2]), 
                .ENAWREN (WREN), 
                .ENBRDEN (RDEN), 
                .REGCEA (REGCE), 
                .REGCEBREGCE (REGCE), 
                .RSTA (1'b0), 
                .RSTBRST (RST), 
                .WEAWEL (WE_PATTERN[1:0]), 
                .WEBWEU (WE_PATTERN[3:2])
                );
            end
            else if (BRAM_SIZE == "18Kb") begin : bram18_sdp_stan
             RAMB16BWER # ( 
                .DOA_REG (DO_REG),
                .DOB_REG (DO_REG),
                .INITP_00 (INITP_00),
                .INITP_01 (INITP_01),
                .INITP_02 (INITP_02), 
                .INITP_03 (INITP_03),
                .INITP_04 (INITP_04),
                .INITP_05 (INITP_05),
                .INITP_06 (INITP_06),
                .INITP_07 (INITP_07),
                .INIT_00 (INIT_00), 
                .INIT_01 (INIT_01),
                .INIT_02 (INIT_02),
                .INIT_03 (INIT_03),
                .INIT_04 (INIT_04),
                .INIT_05 (INIT_05),
                .INIT_06 (INIT_06),
                .INIT_07 (INIT_07),
                .INIT_08 (INIT_08),
                .INIT_09 (INIT_09),
                .INIT_0A (INIT_0A),
                .INIT_0B (INIT_0B),
                .INIT_0C (INIT_0C),
                .INIT_0D (INIT_0D),
                .INIT_0E (INIT_0E),
                .INIT_0F (INIT_0F),
                .INIT_10 (INIT_10),
                .INIT_11 (INIT_11),
                .INIT_12 (INIT_12),
                .INIT_13 (INIT_13),
                .INIT_14 (INIT_14),
                .INIT_15 (INIT_15),
                .INIT_16 (INIT_16),
                .INIT_17 (INIT_17),
                .INIT_18 (INIT_18),
                .INIT_19 (INIT_19),
                .INIT_1A (INIT_1A),
                .INIT_1B (INIT_1B),
                .INIT_1C (INIT_1C),
                .INIT_1D (INIT_1D),
                .INIT_1E (INIT_1E),
                .INIT_1F (INIT_1F),
                .INIT_20 (INIT_20),
                .INIT_21 (INIT_21),
                .INIT_22 (INIT_22),
                .INIT_23 (INIT_23),
                .INIT_24 (INIT_24),
                .INIT_25 (INIT_25),
                .INIT_26 (INIT_26),
                .INIT_27 (INIT_27),
                .INIT_28 (INIT_28),
                .INIT_29 (INIT_29),
                .INIT_2A (INIT_2A),
                .INIT_2B (INIT_2B),
                .INIT_2C (INIT_2C),
                .INIT_2D (INIT_2D),
                .INIT_2E (INIT_2E),
                .INIT_2F (INIT_2F),
                .INIT_30 (INIT_30),
                .INIT_31 (INIT_31),
                .INIT_32 (INIT_32),
                .INIT_33 (INIT_33),
                .INIT_34 (INIT_34),
                .INIT_35 (INIT_35),
                .INIT_36 (INIT_36),
                .INIT_37 (INIT_37),
                .INIT_38 (INIT_38),
                .INIT_39 (INIT_39),
                .INIT_3A (INIT_3A),
                .INIT_3B (INIT_3B),
                .INIT_3C (INIT_3C),
                .INIT_3D (INIT_3D),
                .INIT_3E (INIT_3E),
                .INIT_3F (INIT_3F),
                .INIT_A (init_tmp),
                .INIT_B (init_tmp),
		.INIT_FILE (INIT_FILE),
                .DATA_WIDTH_A (wr_width),
                .DATA_WIDTH_B (rd_width),
                .SIM_COLLISION_CHECK (SIM_COLLISION_CHECK),
                .SIM_DEVICE("SPARTAN6"),
                .SRVAL_A (srval_tmp),
                .SRVAL_B (srval_tmp),
                .WRITE_MODE_A (WRITE_MODE),
                .WRITE_MODE_B (WRITE_MODE)
                )  ram16bwe_tdp (
                .DOA (), 
                .DOB (DO_PATTERN), 
                .DOPA (),
                .DOPB (DOP_PATTERN), 
                .ADDRA(WRADDR_PATTERN), 
                .ADDRB(RDADDR_PATTERN), 
                .CLKA (WRCLK), 
                .CLKB (RDCLK), 
                .DIA (DI_PATTERN), 
                .DIB (32'b0), 
                .DIPA (DIP_PATTERN), 
                .DIPB (4'b0), 
                .ENA (WREN), 
                .ENB (RDEN), 
                .REGCEA (1'b0), 
                .REGCEB (REGCE), 
                .RSTA (1'b0), 
                .RSTB (RST), 
                .WEA (WE_PATTERN), 
                .WEB (4'b0)
                );
            end
          end // end generate spartan6
      endcase
    endgenerate  
endmodule



